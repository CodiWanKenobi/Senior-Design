module tb_System_FromFile();

    reg [0:43] in_data;
    reg [0:59] error_mask;
    reg [0:59] modified_data;
    wire [0:43] out_data;
    wire valid;
    
    RS_Top top(in_data, error_mask, out_data, valid);
    
    integer outFile,inFile;

    initial begin
        outFile = $fopen("Output_Data.txt", "w"); //open file for outputting results to
        inFile = $fopen("RS_Input.txt", "r");
        
        while (! $feof(inFile)) begin           //run until reaching end of file
            $fscanf(inFile, "%h", in_data);  //read in a line of the text file
            $fscanf(inFile, "%h", error_mask);  //read in a line of the text file
//            $ferror(inFile,str);
//            $display("%s",str);
            #50
            $fdisplay(outFile, "Input data: %h", in_data);   //write data 
            $fdisplay(outFile, "Error mask: %h", error_mask);   //write data 
            $fdisplay(outFile, "Corrected data: %h", out_data);   //write data 
            if (((in_data == out_data) && valid) || ((in_data != out_data) && (~valid))) begin
                $fdisplay(outFile, "Success\n");   //write data 
            end else begin
                $fdisplay(outFile, "Failure\n");   //write data 
            end
            $fflush(outFile);
            #50;
        end
    end
endmodule

module RS_Top (in, mask, out, valid);
   input  [0:43] in;
   input  [0:59] mask;
   output [0:43] out;
   output valid;
   
   wire [0:59] encoded;
   wire [0:59] masked;
   assign masked = encoded ^ mask;
   RS_Encoder_Optimized enc(in, encoded);
   RS_Decoder dec(masked, out, valid);
endmodule

module RS_Encoder_Optimized ( in, out );
  input [0:43] in;
  output [0:59] out;
  wire   n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439;
  assign out[0] = in[0];
  assign out[1] = in[1];
  assign out[2] = in[2];
  assign out[3] = in[3];
  assign out[4] = in[4];
  assign out[5] = in[5];
  assign out[6] = in[6];
  assign out[7] = in[7];
  assign out[8] = in[8];
  assign out[9] = in[9];
  assign out[10] = in[10];
  assign out[11] = in[11];
  assign out[12] = in[12];
  assign out[13] = in[13];
  assign out[14] = in[14];
  assign out[15] = in[15];
  assign out[16] = in[16];
  assign out[17] = in[17];
  assign out[18] = in[18];
  assign out[19] = in[19];
  assign out[20] = in[20];
  assign out[21] = in[21];
  assign out[22] = in[22];
  assign out[23] = in[23];
  assign out[24] = in[24];
  assign out[25] = in[25];
  assign out[26] = in[26];
  assign out[27] = in[27];
  assign out[28] = in[28];
  assign out[29] = in[29];
  assign out[30] = in[30];
  assign out[31] = in[31];
  assign out[32] = in[32];
  assign out[33] = in[33];
  assign out[34] = in[34];
  assign out[35] = in[35];
  assign out[36] = in[36];
  assign out[37] = in[37];
  assign out[38] = in[38];
  assign out[39] = in[39];
  assign out[40] = in[40];
  assign out[41] = in[41];
  assign out[42] = in[42];
  assign out[43] = in[43];

  BUFX2 U234 ( .A(n248), .Y(n216) );
  BUFX2 U235 ( .A(n260), .Y(n217) );
  BUFX2 U236 ( .A(n280), .Y(n218) );
  BUFX2 U237 ( .A(n382), .Y(n219) );
  BUFX2 U238 ( .A(n396), .Y(n220) );
  BUFX2 U239 ( .A(n426), .Y(n221) );
  BUFX2 U240 ( .A(n298), .Y(n222) );
  BUFX2 U241 ( .A(n367), .Y(n223) );
  BUFX2 U242 ( .A(n282), .Y(n224) );
  BUFX2 U243 ( .A(n337), .Y(n225) );
  BUFX2 U244 ( .A(n289), .Y(n226) );
  BUFX2 U245 ( .A(n432), .Y(n227) );
  BUFX2 U246 ( .A(n263), .Y(n228) );
  BUFX2 U247 ( .A(n267), .Y(n229) );
  BUFX2 U248 ( .A(n325), .Y(n230) );
  BUFX2 U249 ( .A(n410), .Y(n231) );
  BUFX2 U250 ( .A(n276), .Y(n232) );
  BUFX2 U251 ( .A(n319), .Y(n233) );
  BUFX2 U252 ( .A(n368), .Y(n234) );
  BUFX2 U253 ( .A(n372), .Y(n235) );
  BUFX2 U254 ( .A(n322), .Y(n236) );
  BUFX2 U255 ( .A(n427), .Y(n237) );
  INVX1 U256 ( .A(in[23]), .Y(n268) );
  INVX1 U257 ( .A(in[14]), .Y(n424) );
  MUX2X1 U258 ( .B(n424), .A(in[14]), .S(in[38]), .Y(n413) );
  MUX2X1 U259 ( .B(n268), .A(in[23]), .S(n413), .Y(n311) );
  INVX1 U260 ( .A(n311), .Y(n240) );
  INVX1 U261 ( .A(in[31]), .Y(n407) );
  MUX2X1 U262 ( .B(n407), .A(in[31]), .S(in[11]), .Y(n350) );
  INVX1 U263 ( .A(n350), .Y(n238) );
  INVX1 U264 ( .A(in[0]), .Y(n291) );
  MUX2X1 U265 ( .B(n291), .A(in[0]), .S(in[42]), .Y(n313) );
  MUX2X1 U266 ( .B(n238), .A(n350), .S(n313), .Y(n239) );
  MUX2X1 U267 ( .B(n240), .A(n311), .S(n239), .Y(n385) );
  INVX1 U268 ( .A(in[28]), .Y(n315) );
  INVX1 U269 ( .A(in[27]), .Y(n292) );
  AOI22X1 U270 ( .A(in[27]), .B(in[28]), .C(n315), .D(n292), .Y(n427) );
  INVX1 U271 ( .A(n237), .Y(n428) );
  INVX1 U272 ( .A(in[41]), .Y(n394) );
  INVX1 U273 ( .A(in[19]), .Y(n283) );
  AOI22X1 U274 ( .A(in[19]), .B(in[41]), .C(n394), .D(n283), .Y(n289) );
  MUX2X1 U275 ( .B(n428), .A(n237), .S(n226), .Y(n246) );
  INVX1 U276 ( .A(in[7]), .Y(n383) );
  INVX1 U277 ( .A(in[26]), .Y(n330) );
  INVX1 U278 ( .A(in[5]), .Y(n341) );
  INVX1 U279 ( .A(in[12]), .Y(n374) );
  AOI22X1 U280 ( .A(in[12]), .B(in[5]), .C(n341), .D(n374), .Y(n276) );
  MUX2X1 U281 ( .B(n330), .A(in[26]), .S(n232), .Y(n241) );
  MUX2X1 U282 ( .B(n383), .A(in[7]), .S(n241), .Y(n252) );
  INVX1 U283 ( .A(in[2]), .Y(n284) );
  INVX1 U284 ( .A(in[24]), .Y(n257) );
  INVX1 U285 ( .A(in[20]), .Y(n336) );
  MUX2X1 U286 ( .B(n336), .A(in[20]), .S(in[18]), .Y(n258) );
  MUX2X1 U287 ( .B(n257), .A(in[24]), .S(n258), .Y(n242) );
  MUX2X1 U288 ( .B(n284), .A(in[2]), .S(n242), .Y(n274) );
  INVX1 U289 ( .A(in[33]), .Y(n390) );
  INVX1 U290 ( .A(in[8]), .Y(n338) );
  INVX1 U291 ( .A(in[25]), .Y(n279) );
  INVX1 U292 ( .A(in[17]), .Y(n397) );
  INVX1 U293 ( .A(in[32]), .Y(n278) );
  AOI22X1 U294 ( .A(in[32]), .B(in[17]), .C(n397), .D(n278), .Y(n267) );
  MUX2X1 U295 ( .B(n279), .A(in[25]), .S(n229), .Y(n415) );
  MUX2X1 U296 ( .B(n338), .A(in[8]), .S(n415), .Y(n243) );
  MUX2X1 U297 ( .B(n390), .A(in[33]), .S(n243), .Y(n244) );
  FAX1 U298 ( .A(n252), .B(n274), .C(n244), .YS(n245) );
  FAX1 U299 ( .A(n385), .B(n246), .C(n245), .YS(out[59]) );
  INVX1 U300 ( .A(in[30]), .Y(n430) );
  INVX1 U301 ( .A(in[35]), .Y(n423) );
  AOI22X1 U302 ( .A(in[35]), .B(in[2]), .C(n284), .D(n423), .Y(n298) );
  MUX2X1 U303 ( .B(n430), .A(in[30]), .S(n222), .Y(n256) );
  INVX1 U304 ( .A(n256), .Y(n247) );
  INVX1 U305 ( .A(in[40]), .Y(n302) );
  AOI22X1 U306 ( .A(in[33]), .B(in[40]), .C(n302), .D(n390), .Y(n367) );
  MUX2X1 U307 ( .B(n256), .A(n247), .S(n223), .Y(n310) );
  INVX1 U308 ( .A(n310), .Y(n255) );
  MUX2X1 U309 ( .B(n268), .A(in[23]), .S(n226), .Y(n420) );
  INVX1 U310 ( .A(in[13]), .Y(n293) );
  MUX2X1 U311 ( .B(n293), .A(in[13]), .S(n237), .Y(n362) );
  INVX1 U312 ( .A(in[21]), .Y(n317) );
  INVX1 U313 ( .A(in[16]), .Y(n314) );
  INVX1 U314 ( .A(in[37]), .Y(n290) );
  INVX1 U315 ( .A(in[3]), .Y(n406) );
  AOI22X1 U316 ( .A(in[3]), .B(in[8]), .C(n338), .D(n406), .Y(n368) );
  MUX2X1 U317 ( .B(n290), .A(in[37]), .S(n234), .Y(n353) );
  MUX2X1 U318 ( .B(n314), .A(in[16]), .S(n353), .Y(n405) );
  MUX2X1 U319 ( .B(n317), .A(in[21]), .S(n405), .Y(n288) );
  INVX1 U320 ( .A(in[18]), .Y(n249) );
  INVX1 U321 ( .A(in[36]), .Y(n277) );
  AOI22X1 U322 ( .A(in[36]), .B(in[0]), .C(n291), .D(n277), .Y(n248) );
  MUX2X1 U323 ( .B(n249), .A(in[18]), .S(n216), .Y(n250) );
  MUX2X1 U324 ( .B(n257), .A(in[24]), .S(n250), .Y(n251) );
  FAX1 U325 ( .A(n288), .B(n252), .C(n251), .YS(n253) );
  FAX1 U326 ( .A(n420), .B(n362), .C(n253), .YS(n254) );
  MUX2X1 U327 ( .B(n310), .A(n255), .S(n254), .Y(out[48]) );
  INVX1 U328 ( .A(in[9]), .Y(n266) );
  MUX2X1 U329 ( .B(n266), .A(in[9]), .S(n256), .Y(n294) );
  INVX1 U330 ( .A(in[4]), .Y(n335) );
  AOI22X1 U331 ( .A(in[4]), .B(in[26]), .C(n330), .D(n335), .Y(n282) );
  MUX2X1 U332 ( .B(n383), .A(in[7]), .S(n224), .Y(n392) );
  INVX1 U333 ( .A(n392), .Y(n393) );
  AOI22X1 U334 ( .A(n392), .B(in[24]), .C(n257), .D(n393), .Y(n319) );
  INVX1 U335 ( .A(in[39]), .Y(n421) );
  MUX2X1 U336 ( .B(n421), .A(in[39]), .S(n258), .Y(n381) );
  INVX1 U337 ( .A(n381), .Y(n380) );
  AOI22X1 U338 ( .A(n381), .B(in[25]), .C(n279), .D(n380), .Y(n325) );
  INVX1 U339 ( .A(in[1]), .Y(n408) );
  MUX2X1 U340 ( .B(n408), .A(in[1]), .S(in[43]), .Y(n265) );
  INVX1 U341 ( .A(n265), .Y(n259) );
  MUX2X1 U342 ( .B(n265), .A(n259), .S(n350), .Y(n339) );
  XNOR2X1 U343 ( .A(n230), .B(n339), .Y(n306) );
  INVX1 U344 ( .A(in[15]), .Y(n395) );
  AOI22X1 U345 ( .A(in[13]), .B(in[15]), .C(n395), .D(n293), .Y(n263) );
  INVX1 U346 ( .A(n234), .Y(n369) );
  AOI22X1 U347 ( .A(in[5]), .B(in[36]), .C(n277), .D(n341), .Y(n260) );
  MUX2X1 U348 ( .B(n428), .A(n237), .S(n217), .Y(n261) );
  MUX2X1 U349 ( .B(n369), .A(n234), .S(n261), .Y(n262) );
  FAX1 U350 ( .A(n306), .B(n228), .C(n262), .YS(n264) );
  FAX1 U351 ( .A(n294), .B(n233), .C(n264), .YS(out[55]) );
  INVX1 U352 ( .A(n274), .Y(n275) );
  MUX2X1 U353 ( .B(n317), .A(in[21]), .S(n265), .Y(n365) );
  INVX1 U354 ( .A(n365), .Y(n366) );
  INVX1 U355 ( .A(in[6]), .Y(n351) );
  AOI22X1 U356 ( .A(in[9]), .B(in[6]), .C(n351), .D(n266), .Y(n322) );
  MUX2X1 U357 ( .B(n430), .A(in[30]), .S(n236), .Y(n401) );
  MUX2X1 U358 ( .B(n366), .A(n365), .S(n401), .Y(n272) );
  INVX1 U359 ( .A(n353), .Y(n354) );
  MUX2X1 U360 ( .B(n268), .A(in[23]), .S(n229), .Y(n300) );
  MUX2X1 U361 ( .B(n354), .A(n353), .S(n300), .Y(n271) );
  MUX2X1 U362 ( .B(n315), .A(in[28]), .S(n232), .Y(n269) );
  MUX2X1 U363 ( .B(n291), .A(in[0]), .S(n269), .Y(n270) );
  FAX1 U364 ( .A(n272), .B(n271), .C(n270), .YS(n273) );
  MUX2X1 U365 ( .B(n275), .A(n274), .S(n273), .Y(out[46]) );
  INVX1 U366 ( .A(in[10]), .Y(n425) );
  MUX2X1 U367 ( .B(n425), .A(in[10]), .S(n232), .Y(n348) );
  INVX1 U368 ( .A(in[29]), .Y(n324) );
  AOI22X1 U369 ( .A(in[29]), .B(n277), .C(in[36]), .D(n324), .Y(n372) );
  XNOR2X1 U370 ( .A(n348), .B(n235), .Y(n388) );
  MUX2X1 U371 ( .B(n278), .A(in[32]), .S(n388), .Y(n321) );
  MUX2X1 U372 ( .B(n424), .A(in[14]), .S(n321), .Y(n297) );
  AOI22X1 U373 ( .A(in[25]), .B(in[31]), .C(n407), .D(n279), .Y(n280) );
  MUX2X1 U374 ( .B(n302), .A(in[40]), .S(n218), .Y(n281) );
  MUX2X1 U375 ( .B(n292), .A(in[27]), .S(n281), .Y(n286) );
  MUX2X1 U376 ( .B(n283), .A(in[19]), .S(n224), .Y(n364) );
  MUX2X1 U377 ( .B(n284), .A(in[2]), .S(n364), .Y(n285) );
  FAX1 U378 ( .A(n286), .B(n236), .C(n285), .YS(n287) );
  FAX1 U379 ( .A(n297), .B(n288), .C(n287), .YS(out[52]) );
  INVX1 U380 ( .A(in[34]), .Y(n323) );
  MUX2X1 U381 ( .B(in[34]), .A(n323), .S(n392), .Y(n309) );
  XNOR2X1 U382 ( .A(n365), .B(n309), .Y(n438) );
  MUX2X1 U383 ( .B(n290), .A(in[37]), .S(n226), .Y(n416) );
  MUX2X1 U384 ( .B(n291), .A(in[0]), .S(n416), .Y(n295) );
  INVX1 U385 ( .A(in[22]), .Y(n347) );
  AOI22X1 U386 ( .A(in[27]), .B(in[22]), .C(n347), .D(n292), .Y(n337) );
  MUX2X1 U387 ( .B(n293), .A(in[13]), .S(n225), .Y(n328) );
  FAX1 U388 ( .A(n295), .B(n328), .C(n294), .YS(n296) );
  FAX1 U389 ( .A(n438), .B(n297), .C(n296), .YS(out[57]) );
  INVX1 U390 ( .A(n309), .Y(n308) );
  INVX1 U391 ( .A(n235), .Y(n371) );
  MUX2X1 U392 ( .B(n235), .A(n371), .S(n222), .Y(n345) );
  MUX2X1 U393 ( .B(n351), .A(in[6]), .S(n345), .Y(n299) );
  MUX2X1 U394 ( .B(n374), .A(in[12]), .S(n299), .Y(n305) );
  MUX2X1 U395 ( .B(n395), .A(in[15]), .S(n300), .Y(n301) );
  MUX2X1 U396 ( .B(n302), .A(in[40]), .S(n301), .Y(n303) );
  MUX2X1 U397 ( .B(n347), .A(in[22]), .S(n303), .Y(n304) );
  FAX1 U398 ( .A(n306), .B(n305), .C(n304), .YS(n307) );
  MUX2X1 U399 ( .B(n309), .A(n308), .S(n307), .Y(out[51]) );
  INVX1 U400 ( .A(in[43]), .Y(n312) );
  XNOR2X1 U401 ( .A(n311), .B(n310), .Y(n359) );
  MUX2X1 U402 ( .B(n312), .A(in[43]), .S(n359), .Y(n333) );
  MUX2X1 U403 ( .B(n395), .A(in[15]), .S(n313), .Y(n326) );
  MUX2X1 U404 ( .B(n314), .A(in[16]), .S(n326), .Y(n435) );
  MUX2X1 U405 ( .B(n315), .A(in[28]), .S(n381), .Y(n316) );
  MUX2X1 U406 ( .B(n317), .A(in[21]), .S(n316), .Y(n318) );
  FAX1 U407 ( .A(n435), .B(n233), .C(n318), .YS(n320) );
  FAX1 U408 ( .A(n321), .B(n333), .C(n320), .YS(out[50]) );
  INVX1 U409 ( .A(n333), .Y(n334) );
  MUX2X1 U410 ( .B(n323), .A(in[34]), .S(n236), .Y(n361) );
  MUX2X1 U411 ( .B(n324), .A(in[29]), .S(n361), .Y(n418) );
  INVX1 U412 ( .A(n326), .Y(n327) );
  MUX2X1 U413 ( .B(n327), .A(n326), .S(n230), .Y(n378) );
  MUX2X1 U414 ( .B(n394), .A(in[41]), .S(n328), .Y(n329) );
  MUX2X1 U415 ( .B(n330), .A(in[26]), .S(n329), .Y(n331) );
  FAX1 U416 ( .A(n418), .B(n378), .C(n331), .YS(n332) );
  MUX2X1 U417 ( .B(n334), .A(n333), .S(n332), .Y(out[47]) );
  INVX1 U418 ( .A(n345), .Y(n346) );
  INVX1 U419 ( .A(n435), .Y(n436) );
  AOI22X1 U420 ( .A(in[4]), .B(in[20]), .C(n336), .D(n335), .Y(n410) );
  MUX2X1 U421 ( .B(n436), .A(n435), .S(n231), .Y(n357) );
  MUX2X1 U422 ( .B(n338), .A(in[8]), .S(n225), .Y(n343) );
  MUX2X1 U423 ( .B(in[17]), .A(n397), .S(n339), .Y(n340) );
  MUX2X1 U424 ( .B(n341), .A(in[5]), .S(n340), .Y(n342) );
  FAX1 U425 ( .A(n357), .B(n343), .C(n342), .YS(n344) );
  MUX2X1 U426 ( .B(n346), .A(n345), .S(n344), .Y(out[45]) );
  INVX1 U427 ( .A(n359), .Y(n360) );
  INVX1 U428 ( .A(n348), .Y(n349) );
  MUX2X1 U429 ( .B(n347), .A(in[22]), .S(n362), .Y(n412) );
  MUX2X1 U430 ( .B(n349), .A(n348), .S(n412), .Y(n404) );
  MUX2X1 U431 ( .B(n351), .A(in[6]), .S(n350), .Y(n352) );
  MUX2X1 U432 ( .B(n354), .A(n353), .S(n352), .Y(n355) );
  MUX2X1 U433 ( .B(n408), .A(in[1]), .S(n355), .Y(n356) );
  FAX1 U434 ( .A(n404), .B(n357), .C(n356), .YS(n358) );
  MUX2X1 U435 ( .B(n360), .A(n359), .S(n358), .Y(out[58]) );
  INVX1 U436 ( .A(n378), .Y(n379) );
  INVX1 U437 ( .A(n362), .Y(n363) );
  MUX2X1 U438 ( .B(n363), .A(n362), .S(n361), .Y(n386) );
  MUX2X1 U439 ( .B(n366), .A(n365), .S(n364), .Y(n376) );
  MUX2X1 U440 ( .B(n369), .A(n234), .S(n223), .Y(n370) );
  MUX2X1 U441 ( .B(n235), .A(n371), .S(n370), .Y(n373) );
  MUX2X1 U442 ( .B(n374), .A(in[12]), .S(n373), .Y(n375) );
  FAX1 U443 ( .A(n386), .B(n376), .C(n375), .YS(n377) );
  MUX2X1 U444 ( .B(n379), .A(n378), .S(n377), .Y(out[56]) );
  INVX1 U445 ( .A(n388), .Y(n389) );
  AOI22X1 U446 ( .A(n381), .B(in[17]), .C(n397), .D(n380), .Y(n382) );
  MUX2X1 U447 ( .B(n383), .A(in[7]), .S(n219), .Y(n384) );
  FAX1 U448 ( .A(n386), .B(n385), .C(n384), .YS(n387) );
  MUX2X1 U449 ( .B(n389), .A(n388), .S(n387), .Y(out[54]) );
  MUX2X1 U450 ( .B(n390), .A(in[33]), .S(in[11]), .Y(n391) );
  MUX2X1 U451 ( .B(n393), .A(n392), .S(n391), .Y(n402) );
  INVX1 U452 ( .A(in[38]), .Y(n399) );
  AOI22X1 U453 ( .A(in[41]), .B(in[15]), .C(n395), .D(n394), .Y(n396) );
  MUX2X1 U454 ( .B(n397), .A(in[17]), .S(n220), .Y(n398) );
  MUX2X1 U455 ( .B(n399), .A(in[38]), .S(n398), .Y(n400) );
  FAX1 U456 ( .A(n402), .B(n401), .C(n400), .YS(n403) );
  FAX1 U457 ( .A(n405), .B(n404), .C(n403), .YS(out[53]) );
  INVX1 U458 ( .A(n418), .Y(n419) );
  AOI22X1 U459 ( .A(in[3]), .B(in[31]), .C(n407), .D(n406), .Y(n432) );
  MUX2X1 U460 ( .B(n408), .A(in[1]), .S(in[42]), .Y(n409) );
  FAX1 U461 ( .A(n231), .B(n227), .C(n409), .YS(n411) );
  FAX1 U462 ( .A(n413), .B(n412), .C(n411), .YS(n414) );
  FAX1 U463 ( .A(n416), .B(n415), .C(n414), .YS(n417) );
  MUX2X1 U464 ( .B(n419), .A(n418), .S(n417), .Y(out[49]) );
  INVX1 U465 ( .A(n438), .Y(n439) );
  MUX2X1 U466 ( .B(n421), .A(in[39]), .S(n420), .Y(n422) );
  MUX2X1 U467 ( .B(n423), .A(in[35]), .S(n422), .Y(n433) );
  AOI22X1 U468 ( .A(in[14]), .B(in[10]), .C(n425), .D(n424), .Y(n426) );
  MUX2X1 U469 ( .B(n428), .A(n237), .S(n221), .Y(n429) );
  MUX2X1 U470 ( .B(n430), .A(in[30]), .S(n429), .Y(n431) );
  FAX1 U471 ( .A(n433), .B(n227), .C(n431), .YS(n434) );
  MUX2X1 U472 ( .B(n436), .A(n435), .S(n434), .Y(n437) );
  MUX2X1 U473 ( .B(n439), .A(n438), .S(n437), .Y(out[44]) );
endmodule


module RS_Decoder ( msg, decoded, valid );
  input [0:59] msg;
  output [0:43] decoded;
  output valid;
  wire   \lamb/scale_ts3/genblk1[3].mult/added[1] ,
         \lamb/scale_ts3/genblk1[3].mult/added[2] ,
         \lamb/scale_ts3/genblk1[3].mult/added[3] ,
         \lamb/scale_ts3/genblk1[3].mult/added[4] ,
         \lamb/scale_ts3/genblk1[3].mult/logA[0] ,
         \lamb/scale_ts3/genblk1[3].mult/logA[1] ,
         \lamb/scale_ts3/genblk1[3].mult/logA[2] ,
         \lamb/scale_ts3/genblk1[3].mult/logA[3] ,
         \lamb/scale_ts3/genblk1[2].mult/added[1] ,
         \lamb/scale_ts3/genblk1[2].mult/added[2] ,
         \lamb/scale_ts3/genblk1[2].mult/added[3] ,
         \lamb/scale_ts3/genblk1[2].mult/added[4] ,
         \lamb/scale_ts3/genblk1[2].mult/logA[0] ,
         \lamb/scale_ts3/genblk1[2].mult/logA[1] ,
         \lamb/scale_ts3/genblk1[2].mult/logA[2] ,
         \lamb/scale_ts3/genblk1[2].mult/logA[3] ,
         \lamb/scale_ds3/genblk1[3].mult/added[1] ,
         \lamb/scale_ds3/genblk1[3].mult/added[2] ,
         \lamb/scale_ds3/genblk1[3].mult/added[3] ,
         \lamb/scale_ds3/genblk1[3].mult/added[4] ,
         \lamb/scale_ds3/genblk1[3].mult/logA[0] ,
         \lamb/scale_ds3/genblk1[3].mult/logA[1] ,
         \lamb/scale_ds3/genblk1[3].mult/logA[2] ,
         \lamb/scale_ds3/genblk1[3].mult/logA[3] ,
         \lamb/scale_ds3/genblk1[2].mult/added[1] ,
         \lamb/scale_ds3/genblk1[2].mult/added[2] ,
         \lamb/scale_ds3/genblk1[2].mult/added[3] ,
         \lamb/scale_ds3/genblk1[2].mult/added[4] ,
         \lamb/scale_ds3/genblk1[2].mult/logA[0] ,
         \lamb/scale_ds3/genblk1[2].mult/logA[1] ,
         \lamb/scale_ds3/genblk1[2].mult/logA[2] ,
         \lamb/scale_ds3/genblk1[2].mult/logA[3] ,
         \lamb/scale_bs3/genblk1[1].mult/added[1] ,
         \lamb/scale_bs3/genblk1[1].mult/added[2] ,
         \lamb/scale_bs3/genblk1[1].mult/added[3] ,
         \lamb/scale_bs3/genblk1[1].mult/added[4] ,
         \lamb/scale_bs3/genblk1[1].mult/logA[1] ,
         \lamb/scale_bs3/genblk1[1].mult/logA[2] ,
         \lamb/scale_bs3/genblk1[1].mult/logA[3] ,
         \lamb/scale_bs3/genblk1[0].mult/added[1] ,
         \lamb/scale_bs3/genblk1[0].mult/added[2] ,
         \lamb/scale_bs3/genblk1[0].mult/added[3] ,
         \lamb/scale_bs3/genblk1[0].mult/added[4] ,
         \lamb/scale_bs3/genblk1[0].mult/logB[0] ,
         \lamb/scale_bs3/genblk1[0].mult/logB[1] ,
         \lamb/scale_bs3/genblk1[0].mult/logB[2] ,
         \lamb/scale_bs3/genblk1[0].mult/logB[3] ,
         \lamb/scale_bs3/genblk1[0].mult/logA[0] ,
         \lamb/scale_bs3/genblk1[0].mult/logA[1] ,
         \lamb/scale_bs3/genblk1[0].mult/logA[2] ,
         \lamb/scale_bs3/genblk1[0].mult/logA[3] ,
         \lamb/scale_ls3/genblk1[2].mult/added[1] ,
         \lamb/scale_ls3/genblk1[2].mult/added[2] ,
         \lamb/scale_ls3/genblk1[2].mult/added[3] ,
         \lamb/scale_ls3/genblk1[2].mult/added[4] ,
         \lamb/scale_ls3/genblk1[2].mult/logA[0] ,
         \lamb/scale_ls3/genblk1[2].mult/logA[1] ,
         \lamb/scale_ls3/genblk1[2].mult/logA[2] ,
         \lamb/scale_ls3/genblk1[2].mult/logA[3] ,
         \lamb/scale_ls3/genblk1[1].mult/added[1] ,
         \lamb/scale_ls3/genblk1[1].mult/added[2] ,
         \lamb/scale_ls3/genblk1[1].mult/added[3] ,
         \lamb/scale_ls3/genblk1[1].mult/added[4] ,
         \lamb/scale_ls3/genblk1[1].mult/logA[0] ,
         \lamb/scale_ls3/genblk1[1].mult/logA[2] ,
         \lamb/scale_ls3/genblk1[1].mult/logA[3] ,
         \lamb/scale_ls3/genblk1[0].mult/added[1] ,
         \lamb/scale_ls3/genblk1[0].mult/added[2] ,
         \lamb/scale_ls3/genblk1[0].mult/added[3] ,
         \lamb/scale_ls3/genblk1[0].mult/added[4] ,
         \lamb/scale_ls3/genblk1[0].mult/logB[0] ,
         \lamb/scale_ls3/genblk1[0].mult/logB[1] ,
         \lamb/scale_ls3/genblk1[0].mult/logB[2] ,
         \lamb/scale_ls3/genblk1[0].mult/logB[3] ,
         \lamb/scale_ls3/genblk1[0].mult/logA[0] ,
         \lamb/scale_ls3/genblk1[0].mult/logA[1] ,
         \lamb/scale_ls3/genblk1[0].mult/logA[2] ,
         \lamb/scale_ls3/genblk1[0].mult/logA[3] ,
         \lamb/scale_ts2/genblk1[3].mult/added[1] ,
         \lamb/scale_ts2/genblk1[3].mult/added[2] ,
         \lamb/scale_ts2/genblk1[3].mult/added[3] ,
         \lamb/scale_ts2/genblk1[3].mult/added[4] ,
         \lamb/scale_ts2/genblk1[3].mult/logA[0] ,
         \lamb/scale_ts2/genblk1[3].mult/logA[1] ,
         \lamb/scale_ts2/genblk1[3].mult/logA[2] ,
         \lamb/scale_ts2/genblk1[3].mult/logA[3] ,
         \lamb/scale_ts2/genblk1[2].mult/added[1] ,
         \lamb/scale_ts2/genblk1[2].mult/added[2] ,
         \lamb/scale_ts2/genblk1[2].mult/added[3] ,
         \lamb/scale_ts2/genblk1[2].mult/added[4] ,
         \lamb/scale_ts2/genblk1[2].mult/logA[1] ,
         \lamb/scale_ts2/genblk1[2].mult/logA[2] ,
         \lamb/scale_ts2/genblk1[2].mult/logA[3] ,
         \lamb/scale_ts2/genblk1[1].mult/added[1] ,
         \lamb/scale_ts2/genblk1[1].mult/added[2] ,
         \lamb/scale_ts2/genblk1[1].mult/added[3] ,
         \lamb/scale_ts2/genblk1[1].mult/added[4] ,
         \lamb/scale_ts2/genblk1[1].mult/logA[1] ,
         \lamb/scale_ts2/genblk1[1].mult/logA[2] ,
         \lamb/scale_ts2/genblk1[1].mult/logA[3] ,
         \lamb/scale_ds2/genblk1[3].mult/added[1] ,
         \lamb/scale_ds2/genblk1[3].mult/added[2] ,
         \lamb/scale_ds2/genblk1[3].mult/added[3] ,
         \lamb/scale_ds2/genblk1[3].mult/added[4] ,
         \lamb/scale_ds2/genblk1[3].mult/logA[0] ,
         \lamb/scale_ds2/genblk1[3].mult/logA[1] ,
         \lamb/scale_ds2/genblk1[3].mult/logA[3] ,
         \lamb/scale_ds2/genblk1[2].mult/added[1] ,
         \lamb/scale_ds2/genblk1[2].mult/added[2] ,
         \lamb/scale_ds2/genblk1[2].mult/added[3] ,
         \lamb/scale_ds2/genblk1[2].mult/added[4] ,
         \lamb/scale_ds2/genblk1[2].mult/logA[0] ,
         \lamb/scale_ds2/genblk1[2].mult/logA[1] ,
         \lamb/scale_ds2/genblk1[2].mult/logA[3] ,
         \lamb/scale_ds2/genblk1[1].mult/added[1] ,
         \lamb/scale_ds2/genblk1[1].mult/added[2] ,
         \lamb/scale_ds2/genblk1[1].mult/added[3] ,
         \lamb/scale_ds2/genblk1[1].mult/added[4] ,
         \lamb/scale_ds2/genblk1[1].mult/logA[0] ,
         \lamb/scale_ds2/genblk1[1].mult/logA[1] ,
         \lamb/scale_ds2/genblk1[1].mult/logA[3] ,
         \lamb/scale_bs2/genblk1[1].mult/added[1] ,
         \lamb/scale_bs2/genblk1[1].mult/added[2] ,
         \lamb/scale_bs2/genblk1[1].mult/added[3] ,
         \lamb/scale_bs2/genblk1[1].mult/added[4] ,
         \lamb/scale_bs2/genblk1[0].mult/added[1] ,
         \lamb/scale_bs2/genblk1[0].mult/added[2] ,
         \lamb/scale_bs2/genblk1[0].mult/added[3] ,
         \lamb/scale_bs2/genblk1[0].mult/added[4] ,
         \lamb/scale_bs2/genblk1[0].mult/logA[0] ,
         \lamb/scale_bs2/genblk1[0].mult/logA[1] ,
         \lamb/scale_bs2/genblk1[0].mult/logA[2] ,
         \lamb/scale_bs2/genblk1[0].mult/logA[3] ,
         \lamb/scale_ls2/genblk1[2].mult/added[1] ,
         \lamb/scale_ls2/genblk1[2].mult/added[2] ,
         \lamb/scale_ls2/genblk1[2].mult/added[3] ,
         \lamb/scale_ls2/genblk1[2].mult/added[4] ,
         \lamb/scale_ls2/genblk1[1].mult/added[1] ,
         \lamb/scale_ls2/genblk1[1].mult/added[2] ,
         \lamb/scale_ls2/genblk1[1].mult/added[3] ,
         \lamb/scale_ls2/genblk1[1].mult/added[4] ,
         \lamb/scale_ls2/genblk1[1].mult/logA[2] ,
         \lamb/scale_ls2/genblk1[1].mult/logA[3] ,
         \lamb/scale_ls2/genblk1[0].mult/added[1] ,
         \lamb/scale_ls2/genblk1[0].mult/added[2] ,
         \lamb/scale_ls2/genblk1[0].mult/added[3] ,
         \lamb/scale_ls2/genblk1[0].mult/added[4] ,
         \lamb/scale_ls2/genblk1[0].mult/logB[0] ,
         \lamb/scale_ls2/genblk1[0].mult/logB[1] ,
         \lamb/scale_ls2/genblk1[0].mult/logB[2] ,
         \lamb/scale_ls2/genblk1[0].mult/logB[3] ,
         \lamb/scale_ls2/genblk1[0].mult/logA[0] ,
         \lamb/scale_ls2/genblk1[0].mult/logA[1] ,
         \lamb/scale_ls2/genblk1[0].mult/logA[2] ,
         \lamb/scale_ls2/genblk1[0].mult/logA[3] ,
         \lamb/scale_ts1/genblk1[3].mult/added[1] ,
         \lamb/scale_ts1/genblk1[3].mult/added[2] ,
         \lamb/scale_ts1/genblk1[3].mult/added[3] ,
         \lamb/scale_ts1/genblk1[3].mult/added[4] ,
         \lamb/scale_ts1/genblk1[3].mult/logA[0] ,
         \lamb/scale_ts1/genblk1[2].mult/added[1] ,
         \lamb/scale_ts1/genblk1[2].mult/added[2] ,
         \lamb/scale_ts1/genblk1[2].mult/added[3] ,
         \lamb/scale_ts1/genblk1[2].mult/added[4] ,
         \lamb/scale_ts1/genblk1[2].mult/logA[0] ,
         \lamb/scale_ts1/genblk1[2].mult/logA[1] ,
         \lamb/scale_ts1/genblk1[2].mult/logA[2] ,
         \lamb/scale_ts1/genblk1[2].mult/logA[3] ,
         \lamb/scale_ts1/genblk1[1].mult/added[1] ,
         \lamb/scale_ts1/genblk1[1].mult/added[2] ,
         \lamb/scale_ts1/genblk1[1].mult/added[3] ,
         \lamb/scale_ts1/genblk1[1].mult/added[4] ,
         \lamb/scale_ts1/genblk1[1].mult/logA[0] ,
         \lamb/scale_ts1/genblk1[1].mult/logA[1] ,
         \lamb/scale_ts1/genblk1[1].mult/logA[2] ,
         \lamb/scale_ts1/genblk1[1].mult/logA[3] ,
         \lamb/scale_ts1/genblk1[0].mult/added[1] ,
         \lamb/scale_ts1/genblk1[0].mult/added[2] ,
         \lamb/scale_ts1/genblk1[0].mult/added[3] ,
         \lamb/scale_ts1/genblk1[0].mult/added[4] ,
         \lamb/scale_ts1/genblk1[0].mult/logB[0] ,
         \lamb/scale_ts1/genblk1[0].mult/logB[1] ,
         \lamb/scale_ts1/genblk1[0].mult/logB[2] ,
         \lamb/scale_ts1/genblk1[0].mult/logB[3] ,
         \lamb/scale_ts1/genblk1[0].mult/logA[0] ,
         \lamb/scale_ts1/genblk1[0].mult/logA[1] ,
         \lamb/scale_ts1/genblk1[0].mult/logA[2] ,
         \lamb/scale_ts1/genblk1[0].mult/logA[3] ,
         \lamb/scale_ds1/genblk1[3].mult/added[1] ,
         \lamb/scale_ds1/genblk1[3].mult/added[2] ,
         \lamb/scale_ds1/genblk1[3].mult/added[3] ,
         \lamb/scale_ds1/genblk1[3].mult/added[4] ,
         \lamb/scale_ds1/genblk1[3].mult/logA[1] ,
         \lamb/scale_ds1/genblk1[3].mult/logA[3] ,
         \lamb/scale_ds1/genblk1[2].mult/added[1] ,
         \lamb/scale_ds1/genblk1[2].mult/added[2] ,
         \lamb/scale_ds1/genblk1[2].mult/added[3] ,
         \lamb/scale_ds1/genblk1[2].mult/added[4] ,
         \lamb/scale_ds1/genblk1[2].mult/logA[1] ,
         \lamb/scale_ds1/genblk1[2].mult/logA[2] ,
         \lamb/scale_ds1/genblk1[2].mult/logA[3] ,
         \lamb/scale_ds1/genblk1[1].mult/added[1] ,
         \lamb/scale_ds1/genblk1[1].mult/added[2] ,
         \lamb/scale_ds1/genblk1[1].mult/added[3] ,
         \lamb/scale_ds1/genblk1[1].mult/added[4] ,
         \lamb/scale_ds1/genblk1[1].mult/logA[0] ,
         \lamb/scale_ds1/genblk1[1].mult/logA[1] ,
         \lamb/scale_ds1/genblk1[1].mult/logA[3] ,
         \lamb/scale_ls1/genblk1[1].mult/added[2] ,
         \lamb/scale_ls1/genblk1[1].mult/added[3] ,
         \lamb/scale_ts0/genblk1[2].mult/added[1] ,
         \lamb/scale_ts0/genblk1[2].mult/added[2] ,
         \lamb/scale_ts0/genblk1[2].mult/added[3] ,
         \lamb/scale_ts0/genblk1[2].mult/added[4] ,
         \lamb/scale_ts0/genblk1[2].mult/logA[2] ,
         \lamb/scale_ts0/genblk1[1].mult/added[1] ,
         \lamb/scale_ts0/genblk1[1].mult/added[2] ,
         \lamb/scale_ts0/genblk1[1].mult/added[3] ,
         \lamb/scale_ts0/genblk1[1].mult/added[4] ,
         \lamb/scale_ts0/genblk1[1].mult/logA[1] ,
         \lamb/scale_ts0/genblk1[1].mult/logA[2] ,
         \lamb/scale_ts0/genblk1[1].mult/logA[3] ,
         \lamb/scale_ts0/genblk1[0].mult/added[1] ,
         \lamb/scale_ts0/genblk1[0].mult/added[2] ,
         \lamb/scale_ts0/genblk1[0].mult/added[3] ,
         \lamb/scale_ts0/genblk1[0].mult/added[4] ,
         \lamb/scale_ts0/genblk1[0].mult/logA[0] ,
         \lamb/scale_ts0/genblk1[0].mult/logA[1] ,
         \lamb/scale_ts0/genblk1[0].mult/logA[2] ,
         \lamb/scale_ts0/genblk1[0].mult/logA[3] , \add_x_154/n4 ,
         \add_x_154/n3 , \add_x_154/n2 , \add_x_154/n1 , \add_x_153/n4 ,
         \add_x_153/n3 , \add_x_153/n2 , \add_x_153/n1 , \add_x_152/n4 ,
         \add_x_152/n3 , \add_x_152/n2 , \add_x_152/n1 , \add_x_148/n4 ,
         \add_x_148/n3 , \add_x_148/n2 , \add_x_148/n1 , \add_x_147/n4 ,
         \add_x_147/n3 , \add_x_147/n2 , \add_x_147/n1 , \add_x_146/n4 ,
         \add_x_146/n3 , \add_x_146/n2 , \add_x_146/n1 , \add_x_145/n4 ,
         \add_x_145/n3 , \add_x_145/n2 , \add_x_145/n1 , \add_x_144/n4 ,
         \add_x_144/n3 , \add_x_144/n2 , \add_x_144/n1 , \add_x_143/n4 ,
         \add_x_143/n3 , \add_x_143/n2 , \add_x_143/n1 , \add_x_142/n4 ,
         \add_x_142/n3 , \add_x_142/n2 , \add_x_142/n1 , \add_x_141/n4 ,
         \add_x_141/n3 , \add_x_141/n2 , \add_x_141/n1 , \add_x_140/n4 ,
         \add_x_140/n3 , \add_x_140/n2 , \add_x_140/n1 , \add_x_139/n4 ,
         \add_x_139/n3 , \add_x_139/n2 , \add_x_139/n1 , \add_x_138/n4 ,
         \add_x_138/n3 , \add_x_138/n2 , \add_x_138/n1 , \add_x_135/n4 ,
         \add_x_135/n3 , \add_x_135/n2 , \add_x_135/n1 , \add_x_134/n4 ,
         \add_x_134/n3 , \add_x_134/n2 , \add_x_134/n1 , \add_x_133/n4 ,
         \add_x_133/n3 , \add_x_133/n2 , \add_x_133/n1 , \add_x_131/n4 ,
         \add_x_131/n3 , \add_x_131/n2 , \add_x_131/n1 , \add_x_130/n4 ,
         \add_x_130/n3 , \add_x_130/n2 , \add_x_130/n1 , \add_x_129/n4 ,
         \add_x_129/n3 , \add_x_129/n2 , \add_x_129/n1 , \add_x_128/n4 ,
         \add_x_128/n3 , \add_x_128/n2 , \add_x_128/n1 , \add_x_127/n4 ,
         \add_x_127/n3 , \add_x_127/n2 , \add_x_127/n1 , \add_x_126/n4 ,
         \add_x_126/n3 , \add_x_126/n2 , \add_x_126/n1 , \add_x_125/n4 ,
         \add_x_125/n3 , \add_x_125/n2 , \add_x_125/n1 , \add_x_124/n4 ,
         \add_x_124/n3 , \add_x_124/n2 , \add_x_124/n1 , \add_x_121/n4 ,
         \add_x_121/n3 , \add_x_121/n2 , \add_x_121/n1 , \add_x_120/n4 ,
         \add_x_120/n3 , \add_x_120/n2 , \add_x_120/n1 , \add_x_117/n4 ,
         \add_x_117/n3 , \add_x_117/n2 , \add_x_117/n1 , \add_x_116/n4 ,
         \add_x_116/n3 , \add_x_116/n2 , \add_x_116/n1 , \add_x_87/n4 ,
         \add_x_87/n3 , \add_x_87/n2 , \add_x_87/n1 , \add_x_85/n4 ,
         \add_x_85/n3 , \add_x_85/n2 , \add_x_85/n1 , \add_x_20/n4 ,
         \add_x_20/n3 , \add_x_20/n2 , \add_x_20/n1 , \add_x_14/n4 ,
         \add_x_14/n3 , \add_x_14/n2 , \add_x_14/n1 , n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946;
  wire   [0:4] \forney/m0/added ;
  wire   [0:3] \forney/m0/logB ;
  wire   [0:3] \forney/m0/logA ;
  wire   [0:4] \forney/m1/added ;
  wire   [0:3] \forney/m1/logB ;
  wire   [0:3] \forney/m1/logA ;
  wire   [0:4] \forney/pe1/mult0/added ;
  wire   [0:3] \forney/pe1/mult0/logB ;
  wire   [0:4] \forney/pe0/mult0/added ;
  wire   [0:3] \forney/pe0/mult0/logB ;
  wire   [0:3] \forney/pe0/mult0/logA ;

  HAX1 \add_x_154/U5  ( .A(\lamb/scale_ls1/genblk1[1].mult/added[3] ), .B(
        n10411), .YC(\add_x_154/n4 ), .YS(
        \lamb/scale_ts0/genblk1[0].mult/added[4] ) );
  FAX1 \add_x_154/U4  ( .A(\lamb/scale_ls1/genblk1[1].mult/added[2] ), .B(
        n10786), .C(\add_x_154/n4 ), .YC(\add_x_154/n3 ), .YS(
        \lamb/scale_ts0/genblk1[0].mult/added[3] ) );
  FAX1 \add_x_154/U3  ( .A(n11231), .B(n10787), .C(\add_x_154/n3 ), .YC(
        \add_x_154/n2 ), .YS(\lamb/scale_ts0/genblk1[0].mult/added[2] ) );
  FAX1 \add_x_154/U2  ( .A(n10376), .B(
        \lamb/scale_ts0/genblk1[0].mult/logA[0] ), .C(\add_x_154/n2 ), .YC(
        \add_x_154/n1 ), .YS(\lamb/scale_ts0/genblk1[0].mult/added[1] ) );
  HAX1 \add_x_153/U5  ( .A(\lamb/scale_ls1/genblk1[1].mult/added[3] ), .B(
        \lamb/scale_ts0/genblk1[1].mult/logA[3] ), .YC(\add_x_153/n4 ), .YS(
        \lamb/scale_ts0/genblk1[1].mult/added[4] ) );
  FAX1 \add_x_153/U4  ( .A(\lamb/scale_ls1/genblk1[1].mult/added[2] ), .B(
        n11047), .C(\add_x_153/n4 ), .YC(\add_x_153/n3 ), .YS(
        \lamb/scale_ts0/genblk1[1].mult/added[3] ) );
  FAX1 \add_x_153/U3  ( .A(n11231), .B(n10774), .C(\add_x_153/n3 ), .YC(
        \add_x_153/n2 ), .YS(\lamb/scale_ts0/genblk1[1].mult/added[2] ) );
  FAX1 \add_x_153/U2  ( .A(n10376), .B(n10380), .C(\add_x_153/n2 ), .YC(
        \add_x_153/n1 ), .YS(\lamb/scale_ts0/genblk1[1].mult/added[1] ) );
  HAX1 \add_x_152/U5  ( .A(\lamb/scale_ls1/genblk1[1].mult/added[3] ), .B(
        n10701), .YC(\add_x_152/n4 ), .YS(
        \lamb/scale_ts0/genblk1[2].mult/added[4] ) );
  FAX1 \add_x_152/U4  ( .A(\lamb/scale_ls1/genblk1[1].mult/added[2] ), .B(
        \lamb/scale_ts0/genblk1[2].mult/logA[2] ), .C(\add_x_152/n4 ), .YC(
        \add_x_152/n3 ), .YS(\lamb/scale_ts0/genblk1[2].mult/added[3] ) );
  FAX1 \add_x_152/U3  ( .A(n11231), .B(n10792), .C(\add_x_152/n3 ), .YC(
        \add_x_152/n2 ), .YS(\lamb/scale_ts0/genblk1[2].mult/added[2] ) );
  FAX1 \add_x_152/U2  ( .A(n10376), .B(n10379), .C(\add_x_152/n2 ), .YC(
        \add_x_152/n1 ), .YS(\lamb/scale_ts0/genblk1[2].mult/added[1] ) );
  HAX1 \add_x_148/U5  ( .A(\lamb/scale_ls1/genblk1[1].mult/added[3] ), .B(
        \lamb/scale_ds1/genblk1[1].mult/logA[3] ), .YC(\add_x_148/n4 ), .YS(
        \lamb/scale_ds1/genblk1[1].mult/added[4] ) );
  FAX1 \add_x_148/U4  ( .A(\lamb/scale_ls1/genblk1[1].mult/added[2] ), .B(
        n10362), .C(\add_x_148/n4 ), .YC(\add_x_148/n3 ), .YS(
        \lamb/scale_ds1/genblk1[1].mult/added[3] ) );
  FAX1 \add_x_148/U3  ( .A(n11231), .B(
        \lamb/scale_ds1/genblk1[1].mult/logA[1] ), .C(\add_x_148/n3 ), .YC(
        \add_x_148/n2 ), .YS(\lamb/scale_ds1/genblk1[1].mult/added[2] ) );
  FAX1 \add_x_148/U2  ( .A(n10376), .B(
        \lamb/scale_ds1/genblk1[1].mult/logA[0] ), .C(\add_x_148/n2 ), .YC(
        \add_x_148/n1 ), .YS(\lamb/scale_ds1/genblk1[1].mult/added[1] ) );
  HAX1 \add_x_147/U5  ( .A(\lamb/scale_ls1/genblk1[1].mult/added[3] ), .B(
        \lamb/scale_ds1/genblk1[2].mult/logA[3] ), .YC(\add_x_147/n4 ), .YS(
        \lamb/scale_ds1/genblk1[2].mult/added[4] ) );
  FAX1 \add_x_147/U4  ( .A(\lamb/scale_ls1/genblk1[1].mult/added[2] ), .B(
        n10773), .C(\add_x_147/n4 ), .YC(\add_x_147/n3 ), .YS(
        \lamb/scale_ds1/genblk1[2].mult/added[3] ) );
  FAX1 \add_x_147/U3  ( .A(n11231), .B(
        \lamb/scale_ds1/genblk1[2].mult/logA[1] ), .C(\add_x_147/n3 ), .YC(
        \add_x_147/n2 ), .YS(\lamb/scale_ds1/genblk1[2].mult/added[2] ) );
  FAX1 \add_x_147/U2  ( .A(n10376), .B(n10367), .C(\add_x_147/n2 ), .YC(
        \add_x_147/n1 ), .YS(\lamb/scale_ds1/genblk1[2].mult/added[1] ) );
  HAX1 \add_x_146/U5  ( .A(\lamb/scale_ls1/genblk1[1].mult/added[3] ), .B(
        \lamb/scale_ds1/genblk1[3].mult/logA[3] ), .YC(\add_x_146/n4 ), .YS(
        \lamb/scale_ds1/genblk1[3].mult/added[4] ) );
  FAX1 \add_x_146/U4  ( .A(\lamb/scale_ls1/genblk1[1].mult/added[2] ), .B(
        n10775), .C(\add_x_146/n4 ), .YC(\add_x_146/n3 ), .YS(
        \lamb/scale_ds1/genblk1[3].mult/added[3] ) );
  FAX1 \add_x_146/U3  ( .A(n11231), .B(n10772), .C(\add_x_146/n3 ), .YC(
        \add_x_146/n2 ), .YS(\lamb/scale_ds1/genblk1[3].mult/added[2] ) );
  FAX1 \add_x_146/U2  ( .A(n10376), .B(n10374), .C(\add_x_146/n2 ), .YC(
        \add_x_146/n1 ), .YS(\lamb/scale_ds1/genblk1[3].mult/added[1] ) );
  HAX1 \add_x_145/U5  ( .A(n11206), .B(
        \lamb/scale_ts1/genblk1[0].mult/logA[3] ), .YC(\add_x_145/n4 ), .YS(
        \lamb/scale_ts1/genblk1[0].mult/added[4] ) );
  FAX1 \add_x_145/U4  ( .A(n11214), .B(
        \lamb/scale_ts1/genblk1[0].mult/logA[2] ), .C(\add_x_145/n4 ), .YC(
        \add_x_145/n3 ), .YS(\lamb/scale_ts1/genblk1[0].mult/added[3] ) );
  FAX1 \add_x_145/U3  ( .A(n11213), .B(
        \lamb/scale_ts1/genblk1[0].mult/logA[1] ), .C(\add_x_145/n3 ), .YC(
        \add_x_145/n2 ), .YS(\lamb/scale_ts1/genblk1[0].mult/added[2] ) );
  FAX1 \add_x_145/U2  ( .A(\lamb/scale_ts1/genblk1[0].mult/logB[0] ), .B(
        \lamb/scale_ts1/genblk1[0].mult/logA[0] ), .C(\add_x_145/n2 ), .YC(
        \add_x_145/n1 ), .YS(\lamb/scale_ts1/genblk1[0].mult/added[1] ) );
  HAX1 \add_x_144/U5  ( .A(n11206), .B(
        \lamb/scale_ts1/genblk1[1].mult/logA[3] ), .YC(\add_x_144/n4 ), .YS(
        \lamb/scale_ts1/genblk1[1].mult/added[4] ) );
  FAX1 \add_x_144/U4  ( .A(n11214), .B(n10771), .C(\add_x_144/n4 ), .YC(
        \add_x_144/n3 ), .YS(\lamb/scale_ts1/genblk1[1].mult/added[3] ) );
  FAX1 \add_x_144/U3  ( .A(n11213), .B(
        \lamb/scale_ts1/genblk1[1].mult/logA[1] ), .C(\add_x_144/n3 ), .YC(
        \add_x_144/n2 ), .YS(\lamb/scale_ts1/genblk1[1].mult/added[2] ) );
  FAX1 \add_x_144/U2  ( .A(\lamb/scale_ts1/genblk1[0].mult/logB[0] ), .B(
        \lamb/scale_ts1/genblk1[1].mult/logA[0] ), .C(\add_x_144/n2 ), .YC(
        \add_x_144/n1 ), .YS(\lamb/scale_ts1/genblk1[1].mult/added[1] ) );
  HAX1 \add_x_143/U5  ( .A(n11206), .B(
        \lamb/scale_ts1/genblk1[2].mult/logA[3] ), .YC(\add_x_143/n4 ), .YS(
        \lamb/scale_ts1/genblk1[2].mult/added[4] ) );
  FAX1 \add_x_143/U4  ( .A(n11214), .B(n10770), .C(\add_x_143/n4 ), .YC(
        \add_x_143/n3 ), .YS(\lamb/scale_ts1/genblk1[2].mult/added[3] ) );
  FAX1 \add_x_143/U3  ( .A(n11213), .B(n10769), .C(\add_x_143/n3 ), .YC(
        \add_x_143/n2 ), .YS(\lamb/scale_ts1/genblk1[2].mult/added[2] ) );
  FAX1 \add_x_143/U2  ( .A(\lamb/scale_ts1/genblk1[0].mult/logB[0] ), .B(
        \lamb/scale_ts1/genblk1[2].mult/logA[0] ), .C(\add_x_143/n2 ), .YC(
        \add_x_143/n1 ), .YS(\lamb/scale_ts1/genblk1[2].mult/added[1] ) );
  HAX1 \add_x_142/U5  ( .A(n11206), .B(
        \lamb/scale_ls2/genblk1[1].mult/logA[3] ), .YC(\add_x_142/n4 ), .YS(
        \lamb/scale_ts1/genblk1[3].mult/added[4] ) );
  FAX1 \add_x_142/U4  ( .A(n11214), .B(
        \lamb/scale_ls2/genblk1[1].mult/logA[2] ), .C(\add_x_142/n4 ), .YC(
        \add_x_142/n3 ), .YS(\lamb/scale_ts1/genblk1[3].mult/added[3] ) );
  FAX1 \add_x_142/U3  ( .A(n11213), .B(n10372), .C(\add_x_142/n3 ), .YC(
        \add_x_142/n2 ), .YS(\lamb/scale_ts1/genblk1[3].mult/added[2] ) );
  FAX1 \add_x_142/U2  ( .A(\lamb/scale_ts1/genblk1[0].mult/logB[0] ), .B(
        \lamb/scale_ts1/genblk1[3].mult/logA[0] ), .C(\add_x_142/n2 ), .YC(
        \add_x_142/n1 ), .YS(\lamb/scale_ts1/genblk1[3].mult/added[1] ) );
  HAX1 \add_x_141/U5  ( .A(n10841), .B(
        \lamb/scale_ls2/genblk1[0].mult/logA[3] ), .YC(\add_x_141/n4 ), .YS(
        \lamb/scale_ls2/genblk1[0].mult/added[4] ) );
  FAX1 \add_x_141/U4  ( .A(n11230), .B(
        \lamb/scale_ls2/genblk1[0].mult/logA[2] ), .C(\add_x_141/n4 ), .YC(
        \add_x_141/n3 ), .YS(\lamb/scale_ls2/genblk1[0].mult/added[3] ) );
  FAX1 \add_x_141/U3  ( .A(n10850), .B(
        \lamb/scale_ls2/genblk1[0].mult/logA[1] ), .C(\add_x_141/n3 ), .YC(
        \add_x_141/n2 ), .YS(\lamb/scale_ls2/genblk1[0].mult/added[2] ) );
  FAX1 \add_x_141/U2  ( .A(\lamb/scale_ls2/genblk1[0].mult/logB[0] ), .B(
        \lamb/scale_ls2/genblk1[0].mult/logA[0] ), .C(\add_x_141/n2 ), .YC(
        \add_x_141/n1 ), .YS(\lamb/scale_ls2/genblk1[0].mult/added[1] ) );
  HAX1 \add_x_140/U5  ( .A(n10841), .B(
        \lamb/scale_ls2/genblk1[1].mult/logA[3] ), .YC(\add_x_140/n4 ), .YS(
        \lamb/scale_ls2/genblk1[1].mult/added[4] ) );
  FAX1 \add_x_140/U4  ( .A(n11230), .B(
        \lamb/scale_ls2/genblk1[1].mult/logA[2] ), .C(\add_x_140/n4 ), .YC(
        \add_x_140/n3 ), .YS(\lamb/scale_ls2/genblk1[1].mult/added[3] ) );
  FAX1 \add_x_140/U3  ( .A(n10850), .B(n10372), .C(\add_x_140/n3 ), .YC(
        \add_x_140/n2 ), .YS(\lamb/scale_ls2/genblk1[1].mult/added[2] ) );
  FAX1 \add_x_140/U2  ( .A(\lamb/scale_ls2/genblk1[0].mult/logB[0] ), .B(
        \lamb/scale_ts1/genblk1[3].mult/logA[0] ), .C(\add_x_140/n2 ), .YC(
        \add_x_140/n1 ), .YS(\lamb/scale_ls2/genblk1[1].mult/added[1] ) );
  HAX1 \add_x_139/U5  ( .A(n10841), .B(
        \lamb/scale_ls1/genblk1[1].mult/added[3] ), .YC(\add_x_139/n4 ), .YS(
        \lamb/scale_ls2/genblk1[2].mult/added[4] ) );
  FAX1 \add_x_139/U4  ( .A(n11230), .B(
        \lamb/scale_ls1/genblk1[1].mult/added[2] ), .C(\add_x_139/n4 ), .YC(
        \add_x_139/n3 ), .YS(\lamb/scale_ls2/genblk1[2].mult/added[3] ) );
  FAX1 \add_x_139/U3  ( .A(n10850), .B(n11231), .C(\add_x_139/n3 ), .YC(
        \add_x_139/n2 ), .YS(\lamb/scale_ls2/genblk1[2].mult/added[2] ) );
  FAX1 \add_x_139/U2  ( .A(\lamb/scale_ls2/genblk1[0].mult/logB[0] ), .B(
        n10376), .C(\add_x_139/n2 ), .YC(\add_x_139/n1 ), .YS(
        \lamb/scale_ls2/genblk1[2].mult/added[1] ) );
  HAX1 \add_x_138/U5  ( .A(n11205), .B(
        \lamb/scale_bs2/genblk1[0].mult/logA[3] ), .YC(\add_x_138/n4 ), .YS(
        \lamb/scale_bs2/genblk1[0].mult/added[4] ) );
  FAX1 \add_x_138/U4  ( .A(\lamb/scale_bs2/genblk1[1].mult/added[3] ), .B(
        n10768), .C(\add_x_138/n4 ), .YC(\add_x_138/n3 ), .YS(
        \lamb/scale_bs2/genblk1[0].mult/added[3] ) );
  FAX1 \add_x_138/U3  ( .A(n11212), .B(
        \lamb/scale_bs2/genblk1[0].mult/logA[1] ), .C(\add_x_138/n3 ), .YC(
        \add_x_138/n2 ), .YS(\lamb/scale_bs2/genblk1[0].mult/added[2] ) );
  FAX1 \add_x_138/U2  ( .A(\lamb/scale_bs2/genblk1[1].mult/added[1] ), .B(
        \lamb/scale_bs2/genblk1[0].mult/logA[0] ), .C(\add_x_138/n2 ), .YC(
        \add_x_138/n1 ), .YS(\lamb/scale_bs2/genblk1[0].mult/added[1] ) );
  HAX1 \add_x_135/U5  ( .A(n10841), .B(
        \lamb/scale_ds2/genblk1[1].mult/logA[3] ), .YC(\add_x_135/n4 ), .YS(
        \lamb/scale_ds2/genblk1[1].mult/added[4] ) );
  FAX1 \add_x_135/U4  ( .A(n11230), .B(n10363), .C(\add_x_135/n4 ), .YC(
        \add_x_135/n3 ), .YS(\lamb/scale_ds2/genblk1[1].mult/added[3] ) );
  FAX1 \add_x_135/U3  ( .A(n10850), .B(n10767), .C(\add_x_135/n3 ), .YC(
        \add_x_135/n2 ), .YS(\lamb/scale_ds2/genblk1[1].mult/added[2] ) );
  FAX1 \add_x_135/U2  ( .A(\lamb/scale_ls2/genblk1[0].mult/logB[0] ), .B(
        \lamb/scale_ds2/genblk1[1].mult/logA[0] ), .C(\add_x_135/n2 ), .YC(
        \add_x_135/n1 ), .YS(\lamb/scale_ds2/genblk1[1].mult/added[1] ) );
  HAX1 \add_x_134/U5  ( .A(n10841), .B(
        \lamb/scale_ds2/genblk1[2].mult/logA[3] ), .YC(\add_x_134/n4 ), .YS(
        \lamb/scale_ds2/genblk1[2].mult/added[4] ) );
  FAX1 \add_x_134/U4  ( .A(n11230), .B(n10757), .C(\add_x_134/n4 ), .YC(
        \add_x_134/n3 ), .YS(\lamb/scale_ds2/genblk1[2].mult/added[3] ) );
  FAX1 \add_x_134/U3  ( .A(n10850), .B(n10766), .C(\add_x_134/n3 ), .YC(
        \add_x_134/n2 ), .YS(\lamb/scale_ds2/genblk1[2].mult/added[2] ) );
  FAX1 \add_x_134/U2  ( .A(\lamb/scale_ls2/genblk1[0].mult/logB[0] ), .B(
        \lamb/scale_ds2/genblk1[2].mult/logA[0] ), .C(\add_x_134/n2 ), .YC(
        \add_x_134/n1 ), .YS(\lamb/scale_ds2/genblk1[2].mult/added[1] ) );
  HAX1 \add_x_133/U5  ( .A(n10841), .B(
        \lamb/scale_ds2/genblk1[3].mult/logA[3] ), .YC(\add_x_133/n4 ), .YS(
        \lamb/scale_ds2/genblk1[3].mult/added[4] ) );
  FAX1 \add_x_133/U4  ( .A(n11230), .B(n10777), .C(\add_x_133/n4 ), .YC(
        \add_x_133/n3 ), .YS(\lamb/scale_ds2/genblk1[3].mult/added[3] ) );
  FAX1 \add_x_133/U3  ( .A(n10850), .B(n10756), .C(\add_x_133/n3 ), .YC(
        \add_x_133/n2 ), .YS(\lamb/scale_ds2/genblk1[3].mult/added[2] ) );
  FAX1 \add_x_133/U2  ( .A(\lamb/scale_ls2/genblk1[0].mult/logB[0] ), .B(
        \lamb/scale_ds2/genblk1[3].mult/logA[0] ), .C(\add_x_133/n2 ), .YC(
        \add_x_133/n1 ), .YS(\lamb/scale_ds2/genblk1[3].mult/added[1] ) );
  HAX1 \add_x_131/U5  ( .A(n11205), .B(
        \lamb/scale_ts2/genblk1[1].mult/logA[3] ), .YC(\add_x_131/n4 ), .YS(
        \lamb/scale_ts2/genblk1[1].mult/added[4] ) );
  FAX1 \add_x_131/U4  ( .A(\lamb/scale_bs2/genblk1[1].mult/added[3] ), .B(
        \lamb/scale_ts2/genblk1[1].mult/logA[2] ), .C(\add_x_131/n4 ), .YC(
        \add_x_131/n3 ), .YS(\lamb/scale_ts2/genblk1[1].mult/added[3] ) );
  FAX1 \add_x_131/U3  ( .A(n11212), .B(n10765), .C(\add_x_131/n3 ), .YC(
        \add_x_131/n2 ), .YS(\lamb/scale_ts2/genblk1[1].mult/added[2] ) );
  FAX1 \add_x_131/U2  ( .A(\lamb/scale_bs2/genblk1[1].mult/added[1] ), .B(
        n10360), .C(\add_x_131/n2 ), .YC(\add_x_131/n1 ), .YS(
        \lamb/scale_ts2/genblk1[1].mult/added[1] ) );
  HAX1 \add_x_130/U5  ( .A(n11205), .B(
        \lamb/scale_ts2/genblk1[2].mult/logA[3] ), .YC(\add_x_130/n4 ), .YS(
        \lamb/scale_ts2/genblk1[2].mult/added[4] ) );
  FAX1 \add_x_130/U4  ( .A(\lamb/scale_bs2/genblk1[1].mult/added[3] ), .B(
        n11046), .C(\add_x_130/n4 ), .YC(\add_x_130/n3 ), .YS(
        \lamb/scale_ts2/genblk1[2].mult/added[3] ) );
  FAX1 \add_x_130/U3  ( .A(n11212), .B(
        \lamb/scale_ts2/genblk1[2].mult/logA[1] ), .C(\add_x_130/n3 ), .YC(
        \add_x_130/n2 ), .YS(\lamb/scale_ts2/genblk1[2].mult/added[2] ) );
  FAX1 \add_x_130/U2  ( .A(\lamb/scale_bs2/genblk1[1].mult/added[1] ), .B(
        n10368), .C(\add_x_130/n2 ), .YC(\add_x_130/n1 ), .YS(
        \lamb/scale_ts2/genblk1[2].mult/added[1] ) );
  HAX1 \add_x_129/U5  ( .A(n11205), .B(
        \lamb/scale_ts2/genblk1[3].mult/logA[3] ), .YC(\add_x_129/n4 ), .YS(
        \lamb/scale_ts2/genblk1[3].mult/added[4] ) );
  FAX1 \add_x_129/U4  ( .A(\lamb/scale_bs2/genblk1[1].mult/added[3] ), .B(
        \lamb/scale_ts2/genblk1[3].mult/logA[2] ), .C(\add_x_129/n4 ), .YC(
        \add_x_129/n3 ), .YS(\lamb/scale_ts2/genblk1[3].mult/added[3] ) );
  FAX1 \add_x_129/U3  ( .A(n11212), .B(n10781), .C(\add_x_129/n3 ), .YC(
        \add_x_129/n2 ), .YS(\lamb/scale_ts2/genblk1[3].mult/added[2] ) );
  FAX1 \add_x_129/U2  ( .A(\lamb/scale_bs2/genblk1[1].mult/added[1] ), .B(
        \lamb/scale_ts2/genblk1[3].mult/logA[0] ), .C(\add_x_129/n2 ), .YC(
        \add_x_129/n1 ), .YS(\lamb/scale_ts2/genblk1[3].mult/added[1] ) );
  HAX1 \add_x_128/U5  ( .A(n10834), .B(
        \lamb/scale_ls3/genblk1[0].mult/logA[3] ), .YC(\add_x_128/n4 ), .YS(
        \lamb/scale_ls3/genblk1[0].mult/added[4] ) );
  FAX1 \add_x_128/U4  ( .A(n11226), .B(
        \lamb/scale_ls3/genblk1[0].mult/logA[2] ), .C(\add_x_128/n4 ), .YC(
        \add_x_128/n3 ), .YS(\lamb/scale_ls3/genblk1[0].mult/added[3] ) );
  FAX1 \add_x_128/U3  ( .A(n10844), .B(n10764), .C(\add_x_128/n3 ), .YC(
        \add_x_128/n2 ), .YS(\lamb/scale_ls3/genblk1[0].mult/added[2] ) );
  FAX1 \add_x_128/U2  ( .A(\lamb/scale_ls3/genblk1[0].mult/logB[0] ), .B(
        n10779), .C(\add_x_128/n2 ), .YC(\add_x_128/n1 ), .YS(
        \lamb/scale_ls3/genblk1[0].mult/added[1] ) );
  HAX1 \add_x_127/U5  ( .A(n10834), .B(
        \lamb/scale_ls3/genblk1[1].mult/logA[3] ), .YC(\add_x_127/n4 ), .YS(
        \lamb/scale_ls3/genblk1[1].mult/added[4] ) );
  FAX1 \add_x_127/U4  ( .A(n11226), .B(n10763), .C(\add_x_127/n4 ), .YC(
        \add_x_127/n3 ), .YS(\lamb/scale_ls3/genblk1[1].mult/added[3] ) );
  FAX1 \add_x_127/U3  ( .A(n10844), .B(n10776), .C(\add_x_127/n3 ), .YC(
        \add_x_127/n2 ), .YS(\lamb/scale_ls3/genblk1[1].mult/added[2] ) );
  FAX1 \add_x_127/U2  ( .A(\lamb/scale_ls3/genblk1[0].mult/logB[0] ), .B(
        \lamb/scale_ls3/genblk1[1].mult/logA[0] ), .C(\add_x_127/n2 ), .YC(
        \add_x_127/n1 ), .YS(\lamb/scale_ls3/genblk1[1].mult/added[1] ) );
  HAX1 \add_x_126/U5  ( .A(n10834), .B(
        \lamb/scale_ls3/genblk1[2].mult/logA[3] ), .YC(\add_x_126/n4 ), .YS(
        \lamb/scale_ls3/genblk1[2].mult/added[4] ) );
  FAX1 \add_x_126/U4  ( .A(n11226), .B(
        \lamb/scale_ls3/genblk1[2].mult/logA[2] ), .C(\add_x_126/n4 ), .YC(
        \add_x_126/n3 ), .YS(\lamb/scale_ls3/genblk1[2].mult/added[3] ) );
  FAX1 \add_x_126/U3  ( .A(n10844), .B(n10780), .C(\add_x_126/n3 ), .YC(
        \add_x_126/n2 ), .YS(\lamb/scale_ls3/genblk1[2].mult/added[2] ) );
  FAX1 \add_x_126/U2  ( .A(\lamb/scale_ls3/genblk1[0].mult/logB[0] ), .B(
        n10762), .C(\add_x_126/n2 ), .YC(\add_x_126/n1 ), .YS(
        \lamb/scale_ls3/genblk1[2].mult/added[1] ) );
  HAX1 \add_x_125/U5  ( .A(n11204), .B(
        \lamb/scale_bs3/genblk1[0].mult/logA[3] ), .YC(\add_x_125/n4 ), .YS(
        \lamb/scale_bs3/genblk1[0].mult/added[4] ) );
  FAX1 \add_x_125/U4  ( .A(\lamb/scale_bs3/genblk1[0].mult/logB[2] ), .B(
        \lamb/scale_bs3/genblk1[0].mult/logA[2] ), .C(\add_x_125/n4 ), .YC(
        \add_x_125/n3 ), .YS(\lamb/scale_bs3/genblk1[0].mult/added[3] ) );
  FAX1 \add_x_125/U3  ( .A(n11211), .B(
        \lamb/scale_bs3/genblk1[0].mult/logA[1] ), .C(\add_x_125/n3 ), .YC(
        \add_x_125/n2 ), .YS(\lamb/scale_bs3/genblk1[0].mult/added[2] ) );
  FAX1 \add_x_125/U2  ( .A(\lamb/scale_bs3/genblk1[0].mult/logB[0] ), .B(
        \lamb/scale_bs3/genblk1[0].mult/logA[0] ), .C(\add_x_125/n2 ), .YC(
        \add_x_125/n1 ), .YS(\lamb/scale_bs3/genblk1[0].mult/added[1] ) );
  HAX1 \add_x_124/U5  ( .A(n11204), .B(
        \lamb/scale_bs3/genblk1[1].mult/logA[3] ), .YC(\add_x_124/n4 ), .YS(
        \lamb/scale_bs3/genblk1[1].mult/added[4] ) );
  FAX1 \add_x_124/U4  ( .A(\lamb/scale_bs3/genblk1[0].mult/logB[2] ), .B(
        \lamb/scale_bs3/genblk1[1].mult/logA[2] ), .C(\add_x_124/n4 ), .YC(
        \add_x_124/n3 ), .YS(\lamb/scale_bs3/genblk1[1].mult/added[3] ) );
  FAX1 \add_x_124/U3  ( .A(n11211), .B(n10778), .C(\add_x_124/n3 ), .YC(
        \add_x_124/n2 ), .YS(\lamb/scale_bs3/genblk1[1].mult/added[2] ) );
  FAX1 \add_x_124/U2  ( .A(\lamb/scale_bs3/genblk1[0].mult/logB[0] ), .B(
        n10370), .C(\add_x_124/n2 ), .YC(\add_x_124/n1 ), .YS(
        \lamb/scale_bs3/genblk1[1].mult/added[1] ) );
  HAX1 \add_x_121/U5  ( .A(n10834), .B(
        \lamb/scale_ds3/genblk1[2].mult/logA[3] ), .YC(\add_x_121/n4 ), .YS(
        \lamb/scale_ds3/genblk1[2].mult/added[4] ) );
  FAX1 \add_x_121/U4  ( .A(n11226), .B(n10761), .C(\add_x_121/n4 ), .YC(
        \add_x_121/n3 ), .YS(\lamb/scale_ds3/genblk1[2].mult/added[3] ) );
  FAX1 \add_x_121/U3  ( .A(n10844), .B(n10760), .C(\add_x_121/n3 ), .YC(
        \add_x_121/n2 ), .YS(\lamb/scale_ds3/genblk1[2].mult/added[2] ) );
  FAX1 \add_x_121/U2  ( .A(\lamb/scale_ls3/genblk1[0].mult/logB[0] ), .B(
        \lamb/scale_ds3/genblk1[2].mult/logA[0] ), .C(\add_x_121/n2 ), .YC(
        \add_x_121/n1 ), .YS(\lamb/scale_ds3/genblk1[2].mult/added[1] ) );
  HAX1 \add_x_120/U5  ( .A(n10834), .B(
        \lamb/scale_ds3/genblk1[3].mult/logA[3] ), .YC(\add_x_120/n4 ), .YS(
        \lamb/scale_ds3/genblk1[3].mult/added[4] ) );
  FAX1 \add_x_120/U4  ( .A(n11226), .B(n10758), .C(\add_x_120/n4 ), .YC(
        \add_x_120/n3 ), .YS(\lamb/scale_ds3/genblk1[3].mult/added[3] ) );
  FAX1 \add_x_120/U3  ( .A(n10844), .B(
        \lamb/scale_ds3/genblk1[3].mult/logA[1] ), .C(\add_x_120/n3 ), .YC(
        \add_x_120/n2 ), .YS(\lamb/scale_ds3/genblk1[3].mult/added[2] ) );
  FAX1 \add_x_120/U2  ( .A(\lamb/scale_ls3/genblk1[0].mult/logB[0] ), .B(
        \lamb/scale_ds3/genblk1[3].mult/logA[0] ), .C(\add_x_120/n2 ), .YC(
        \add_x_120/n1 ), .YS(\lamb/scale_ds3/genblk1[3].mult/added[1] ) );
  HAX1 \add_x_117/U5  ( .A(n11204), .B(
        \lamb/scale_ts3/genblk1[2].mult/logA[3] ), .YC(\add_x_117/n4 ), .YS(
        \lamb/scale_ts3/genblk1[2].mult/added[4] ) );
  FAX1 \add_x_117/U4  ( .A(\lamb/scale_bs3/genblk1[0].mult/logB[2] ), .B(
        n11039), .C(\add_x_117/n4 ), .YC(\add_x_117/n3 ), .YS(
        \lamb/scale_ts3/genblk1[2].mult/added[3] ) );
  FAX1 \add_x_117/U3  ( .A(n11211), .B(
        \lamb/scale_ts3/genblk1[2].mult/logA[1] ), .C(\add_x_117/n3 ), .YC(
        \add_x_117/n2 ), .YS(\lamb/scale_ts3/genblk1[2].mult/added[2] ) );
  FAX1 \add_x_117/U2  ( .A(\lamb/scale_bs3/genblk1[0].mult/logB[0] ), .B(
        \lamb/scale_ts3/genblk1[2].mult/logA[0] ), .C(\add_x_117/n2 ), .YC(
        \add_x_117/n1 ), .YS(\lamb/scale_ts3/genblk1[2].mult/added[1] ) );
  HAX1 \add_x_116/U5  ( .A(n11204), .B(
        \lamb/scale_ts3/genblk1[3].mult/logA[3] ), .YC(\add_x_116/n4 ), .YS(
        \lamb/scale_ts3/genblk1[3].mult/added[4] ) );
  FAX1 \add_x_116/U4  ( .A(\lamb/scale_bs3/genblk1[0].mult/logB[2] ), .B(
        n11033), .C(\add_x_116/n4 ), .YC(\add_x_116/n3 ), .YS(
        \lamb/scale_ts3/genblk1[3].mult/added[3] ) );
  FAX1 \add_x_116/U3  ( .A(n11211), .B(
        \lamb/scale_ts3/genblk1[3].mult/logA[1] ), .C(\add_x_116/n3 ), .YC(
        \add_x_116/n2 ), .YS(\lamb/scale_ts3/genblk1[3].mult/added[2] ) );
  FAX1 \add_x_116/U2  ( .A(\lamb/scale_bs3/genblk1[0].mult/logB[0] ), .B(
        \lamb/scale_ts3/genblk1[3].mult/logA[0] ), .C(\add_x_116/n2 ), .YC(
        \add_x_116/n1 ), .YS(\lamb/scale_ts3/genblk1[3].mult/added[1] ) );
  HAX1 \add_x_87/U5  ( .A(\forney/pe0/mult0/logB [3]), .B(
        \forney/pe0/mult0/logA [3]), .YC(\add_x_87/n4 ), .YS(
        \forney/pe0/mult0/added [4]) );
  FAX1 \add_x_87/U4  ( .A(\forney/pe0/mult0/logB [2]), .B(n11178), .C(
        \add_x_87/n4 ), .YC(\add_x_87/n3 ), .YS(\forney/pe0/mult0/added [3])
         );
  FAX1 \add_x_87/U3  ( .A(n10790), .B(\forney/pe0/mult0/logA [1]), .C(
        \add_x_87/n3 ), .YC(\add_x_87/n2 ), .YS(\forney/pe0/mult0/added [2])
         );
  FAX1 \add_x_87/U2  ( .A(\forney/pe0/mult0/logB [0]), .B(
        \forney/pe0/mult0/logA [0]), .C(\add_x_87/n2 ), .YC(\add_x_87/n1 ), 
        .YS(\forney/pe0/mult0/added [1]) );
  HAX1 \add_x_85/U5  ( .A(\forney/pe1/mult0/logB [3]), .B(
        \forney/pe0/mult0/logA [3]), .YC(\add_x_85/n4 ), .YS(
        \forney/pe1/mult0/added [4]) );
  FAX1 \add_x_85/U4  ( .A(\forney/pe1/mult0/logB [2]), .B(n11178), .C(
        \add_x_85/n4 ), .YC(\add_x_85/n3 ), .YS(\forney/pe1/mult0/added [3])
         );
  FAX1 \add_x_85/U3  ( .A(n10789), .B(\forney/pe0/mult0/logA [1]), .C(
        \add_x_85/n3 ), .YC(\add_x_85/n2 ), .YS(\forney/pe1/mult0/added [2])
         );
  FAX1 \add_x_85/U2  ( .A(\forney/pe1/mult0/logB [0]), .B(
        \forney/pe0/mult0/logA [0]), .C(\add_x_85/n2 ), .YC(\add_x_85/n1 ), 
        .YS(\forney/pe1/mult0/added [1]) );
  HAX1 \add_x_20/U5  ( .A(\forney/m1/logB [3]), .B(\forney/m1/logA [3]), .YC(
        \add_x_20/n4 ), .YS(\forney/m1/added [4]) );
  FAX1 \add_x_20/U4  ( .A(\forney/m1/logB [2]), .B(n11032), .C(\add_x_20/n4 ), 
        .YC(\add_x_20/n3 ), .YS(\forney/m1/added [3]) );
  FAX1 \add_x_20/U3  ( .A(n10788), .B(n10791), .C(\add_x_20/n3 ), .YC(
        \add_x_20/n2 ), .YS(\forney/m1/added [2]) );
  FAX1 \add_x_20/U2  ( .A(\forney/m1/logB [0]), .B(n10785), .C(\add_x_20/n2 ), 
        .YC(\add_x_20/n1 ), .YS(\forney/m1/added [1]) );
  HAX1 \add_x_14/U5  ( .A(n10981), .B(\forney/m0/logA [3]), .YC(\add_x_14/n4 ), 
        .YS(\forney/m0/added [4]) );
  FAX1 \add_x_14/U4  ( .A(\forney/m0/logB [2]), .B(\forney/m0/logA [2]), .C(
        \add_x_14/n4 ), .YC(\add_x_14/n3 ), .YS(\forney/m0/added [3]) );
  FAX1 \add_x_14/U3  ( .A(\forney/m0/logB [1]), .B(\forney/m0/logA [1]), .C(
        \add_x_14/n3 ), .YC(\add_x_14/n2 ), .YS(\forney/m0/added [2]) );
  FAX1 \add_x_14/U2  ( .A(\forney/m0/logB [0]), .B(n10759), .C(\add_x_14/n2 ), 
        .YC(\add_x_14/n1 ), .YS(\forney/m0/added [1]) );
  AND2X1 U6889 ( .A(n13487), .B(n10437), .Y(n13696) );
  AND2X1 U6890 ( .A(n10444), .B(n12691), .Y(n13176) );
  AND2X1 U6891 ( .A(n10851), .B(n10411), .Y(
        \lamb/scale_ts1/genblk1[0].mult/logA[3] ) );
  OR2X1 U6892 ( .A(n13325), .B(n10440), .Y(n13224) );
  BUFX2 U6893 ( .A(n13208), .Y(n10381) );
  AND2X1 U6894 ( .A(n11141), .B(n13408), .Y(n13414) );
  INVX1 U6895 ( .A(n13414), .Y(n10382) );
  BUFX2 U6896 ( .A(n12897), .Y(n10383) );
  AND2X1 U6897 ( .A(n13582), .B(n11198), .Y(n13907) );
  INVX1 U6898 ( .A(n13907), .Y(n10384) );
  BUFX2 U6899 ( .A(n11461), .Y(n10385) );
  BUFX2 U6900 ( .A(n11745), .Y(n10386) );
  BUFX2 U6901 ( .A(n11741), .Y(n10387) );
  BUFX2 U6902 ( .A(n11933), .Y(n10388) );
  AND2X1 U6903 ( .A(n10809), .B(n13850), .Y(n11850) );
  INVX1 U6904 ( .A(n11850), .Y(n10389) );
  AND2X2 U6905 ( .A(n12404), .B(n11155), .Y(n12405) );
  INVX1 U6906 ( .A(n12405), .Y(n10390) );
  AND2X1 U6907 ( .A(n11157), .B(n12873), .Y(n12528) );
  INVX1 U6908 ( .A(n12528), .Y(n10391) );
  AND2X2 U6909 ( .A(n12589), .B(n11146), .Y(n12590) );
  INVX1 U6910 ( .A(n12590), .Y(n10392) );
  AND2X2 U6911 ( .A(n12617), .B(n11146), .Y(n12618) );
  INVX1 U6912 ( .A(n12618), .Y(n10393) );
  BUFX2 U6913 ( .A(n12580), .Y(n10394) );
  BUFX2 U6914 ( .A(n13633), .Y(n10395) );
  AND2X1 U6915 ( .A(n13248), .B(n13249), .Y(n12712) );
  INVX1 U6916 ( .A(n12712), .Y(n10396) );
  AND2X1 U6917 ( .A(\add_x_143/n1 ), .B(
        \lamb/scale_ts1/genblk1[2].mult/added[4] ), .Y(n11639) );
  INVX1 U6918 ( .A(n11639), .Y(n10397) );
  BUFX2 U6919 ( .A(n12919), .Y(n10398) );
  BUFX2 U6920 ( .A(n13103), .Y(n10399) );
  BUFX2 U6921 ( .A(n13197), .Y(n10400) );
  BUFX2 U6922 ( .A(n13277), .Y(n10401) );
  BUFX2 U6923 ( .A(n13125), .Y(n10402) );
  AND2X1 U6924 ( .A(n13934), .B(n13204), .Y(n13939) );
  INVX1 U6925 ( .A(n13939), .Y(n10403) );
  BUFX2 U6926 ( .A(n12927), .Y(n10404) );
  BUFX2 U6927 ( .A(n12575), .Y(n10405) );
  BUFX2 U6928 ( .A(n12472), .Y(n10406) );
  AND2X1 U6929 ( .A(n13937), .B(n13934), .Y(n13940) );
  INVX1 U6930 ( .A(n13940), .Y(n10407) );
  BUFX2 U6931 ( .A(n12413), .Y(n10408) );
  AND2X1 U6932 ( .A(n12858), .B(n12810), .Y(n12815) );
  INVX1 U6933 ( .A(n12815), .Y(n10409) );
  BUFX2 U6934 ( .A(n13621), .Y(n10410) );
  BUFX2 U6935 ( .A(\lamb/scale_ts0/genblk1[0].mult/logA[3] ), .Y(n10411) );
  INVX1 U6936 ( .A(n10412), .Y(n13918) );
  INVX1 U6937 ( .A(n13211), .Y(n10413) );
  INVX1 U6938 ( .A(n10646), .Y(n10414) );
  INVX1 U6939 ( .A(n13222), .Y(n10415) );
  NOR2X1 U6940 ( .A(n10415), .B(n10416), .Y(n10412) );
  NOR2X1 U6941 ( .A(n10413), .B(n10414), .Y(n10417) );
  INVX1 U6942 ( .A(n10417), .Y(n10416) );
  BUFX2 U6943 ( .A(n13611), .Y(n10418) );
  BUFX2 U6944 ( .A(n13642), .Y(n10419) );
  AND2X1 U6945 ( .A(n13318), .B(n13327), .Y(n13330) );
  INVX1 U6946 ( .A(n13330), .Y(n10420) );
  BUFX2 U6947 ( .A(n11807), .Y(n10421) );
  BUFX2 U6948 ( .A(n11752), .Y(n10422) );
  AND2X1 U6949 ( .A(\lamb/scale_ds1/genblk1[3].mult/added[2] ), .B(n11106), 
        .Y(n11424) );
  INVX1 U6950 ( .A(n11424), .Y(n10423) );
  OR2X1 U6951 ( .A(n11075), .B(n10808), .Y(n13283) );
  INVX1 U6952 ( .A(n13283), .Y(n10424) );
  OR2X1 U6953 ( .A(n13868), .B(n12690), .Y(n13173) );
  INVX1 U6954 ( .A(n13173), .Y(n10425) );
  BUFX2 U6955 ( .A(n12903), .Y(n10426) );
  AND2X1 U6956 ( .A(\lamb/scale_ds2/genblk1[3].mult/added[2] ), .B(
        \lamb/scale_ds2/genblk1[3].mult/added[1] ), .Y(n11758) );
  INVX1 U6957 ( .A(n11758), .Y(n10427) );
  AND2X1 U6958 ( .A(\lamb/scale_ts3/genblk1[2].mult/added[1] ), .B(
        \lamb/scale_ts3/genblk1[2].mult/added[2] ), .Y(n12389) );
  INVX1 U6959 ( .A(n12389), .Y(n10428) );
  AND2X1 U6960 ( .A(n11108), .B(n13555), .Y(n13541) );
  INVX1 U6961 ( .A(n13541), .Y(n10429) );
  BUFX2 U6962 ( .A(n13282), .Y(n10430) );
  BUFX2 U6963 ( .A(n13036), .Y(n10431) );
  BUFX2 U6964 ( .A(n13172), .Y(n10432) );
  BUFX2 U6965 ( .A(n12402), .Y(n10433) );
  BUFX2 U6966 ( .A(n12464), .Y(n10434) );
  BUFX2 U6967 ( .A(n12883), .Y(n10435) );
  AND2X1 U6968 ( .A(\lamb/scale_ds3/genblk1[2].mult/added[1] ), .B(n12401), 
        .Y(n12420) );
  INVX1 U6969 ( .A(n12420), .Y(n10436) );
  AND2X1 U6970 ( .A(n12804), .B(n12822), .Y(n12786) );
  INVX1 U6971 ( .A(n12786), .Y(n10437) );
  AND2X1 U6972 ( .A(n10445), .B(n13443), .Y(n13449) );
  INVX1 U6973 ( .A(n13449), .Y(n10438) );
  OR2X1 U6974 ( .A(n12916), .B(n12911), .Y(n13491) );
  INVX1 U6975 ( .A(n13491), .Y(n10439) );
  AND2X1 U6976 ( .A(n13326), .B(n13317), .Y(n13319) );
  INVX1 U6977 ( .A(n13319), .Y(n10440) );
  AND2X1 U6978 ( .A(\lamb/scale_ls3/genblk1[2].mult/added[3] ), .B(n11944), 
        .Y(n11935) );
  INVX1 U6979 ( .A(n11935), .Y(n10441) );
  BUFX2 U6980 ( .A(n12800), .Y(n10442) );
  BUFX2 U6981 ( .A(n11617), .Y(n10443) );
  BUFX2 U6982 ( .A(n12689), .Y(n10444) );
  AND2X2 U6983 ( .A(n11202), .B(n13412), .Y(n13445) );
  INVX1 U6984 ( .A(n13445), .Y(n10445) );
  AND2X2 U6985 ( .A(n12215), .B(n12214), .Y(n12270) );
  AND2X2 U6986 ( .A(n11857), .B(n12304), .Y(n11453) );
  AND2X2 U6987 ( .A(n13903), .B(n12772), .Y(\forney/m0/logA [1]) );
  AND2X2 U6988 ( .A(n12446), .B(n12445), .Y(n12498) );
  AND2X2 U6989 ( .A(n13596), .B(n12824), .Y(n12847) );
  AND2X2 U6990 ( .A(n10830), .B(n13038), .Y(n13041) );
  AND2X2 U6991 ( .A(n13273), .B(n13275), .Y(n13264) );
  INVX1 U6992 ( .A(n10448), .Y(n10446) );
  INVX1 U6993 ( .A(n10446), .Y(n10447) );
  BUFX2 U6994 ( .A(n12850), .Y(n10448) );
  INVX1 U6995 ( .A(n10451), .Y(n10449) );
  INVX1 U6996 ( .A(n10449), .Y(n10450) );
  BUFX2 U6997 ( .A(n12834), .Y(n10451) );
  INVX1 U6998 ( .A(n10454), .Y(n10452) );
  INVX1 U6999 ( .A(n10452), .Y(n10453) );
  OR2X1 U7000 ( .A(n11169), .B(n13248), .Y(n12710) );
  INVX1 U7001 ( .A(n12710), .Y(n10454) );
  INVX1 U7002 ( .A(n10457), .Y(n10455) );
  INVX1 U7003 ( .A(n10455), .Y(n10456) );
  BUFX2 U7004 ( .A(n13530), .Y(n10457) );
  INVX1 U7005 ( .A(n10460), .Y(n10458) );
  INVX1 U7006 ( .A(n10458), .Y(n10459) );
  BUFX2 U7007 ( .A(n13511), .Y(n10460) );
  INVX1 U7008 ( .A(n10463), .Y(n10461) );
  INVX1 U7009 ( .A(n10461), .Y(n10462) );
  AND2X1 U7010 ( .A(n10676), .B(n13841), .Y(n11904) );
  INVX1 U7011 ( .A(n11904), .Y(n10463) );
  INVX1 U7012 ( .A(n10466), .Y(n10464) );
  INVX1 U7013 ( .A(n10464), .Y(n10465) );
  AND2X1 U7014 ( .A(n12682), .B(n10630), .Y(n12366) );
  INVX1 U7015 ( .A(n12366), .Y(n10466) );
  INVX1 U7016 ( .A(n10469), .Y(n10467) );
  INVX1 U7017 ( .A(n10467), .Y(n10468) );
  AND2X1 U7018 ( .A(n12335), .B(n11134), .Y(n13923) );
  INVX1 U7019 ( .A(n13923), .Y(n10469) );
  INVX1 U7020 ( .A(n10472), .Y(n10470) );
  INVX1 U7021 ( .A(n10470), .Y(n10471) );
  BUFX2 U7022 ( .A(n13261), .Y(n10472) );
  INVX1 U7023 ( .A(n10475), .Y(n10473) );
  INVX1 U7024 ( .A(n10473), .Y(n10474) );
  AND2X1 U7025 ( .A(n12335), .B(n13925), .Y(n13361) );
  INVX1 U7026 ( .A(n13361), .Y(n10475) );
  INVX1 U7027 ( .A(n10478), .Y(n10476) );
  INVX1 U7028 ( .A(n10476), .Y(n10477) );
  INVX1 U7029 ( .A(n13696), .Y(n10478) );
  INVX1 U7030 ( .A(n10481), .Y(n10479) );
  INVX1 U7031 ( .A(n10479), .Y(n10480) );
  BUFX2 U7032 ( .A(n13887), .Y(n10481) );
  INVX1 U7033 ( .A(n10484), .Y(n10482) );
  INVX1 U7034 ( .A(n10482), .Y(n10483) );
  BUFX2 U7035 ( .A(n13137), .Y(n10484) );
  INVX1 U7036 ( .A(n10487), .Y(n10485) );
  INVX1 U7037 ( .A(n10485), .Y(n10486) );
  AND2X1 U7038 ( .A(n13100), .B(n13097), .Y(n13090) );
  INVX1 U7039 ( .A(n13090), .Y(n10487) );
  INVX1 U7040 ( .A(n10490), .Y(n10488) );
  INVX1 U7041 ( .A(n10488), .Y(n10489) );
  AND2X1 U7042 ( .A(n13846), .B(n13858), .Y(n13849) );
  INVX1 U7043 ( .A(n13849), .Y(n10490) );
  INVX1 U7044 ( .A(n10493), .Y(n10491) );
  INVX1 U7045 ( .A(n10491), .Y(n10492) );
  INVX1 U7046 ( .A(n13176), .Y(n10493) );
  INVX1 U7047 ( .A(n10496), .Y(n10494) );
  INVX1 U7048 ( .A(n10494), .Y(n10495) );
  AND2X1 U7049 ( .A(n10703), .B(n10800), .Y(n13942) );
  INVX1 U7050 ( .A(n13942), .Y(n10496) );
  INVX1 U7051 ( .A(n10499), .Y(n10497) );
  INVX1 U7052 ( .A(n10497), .Y(n10498) );
  AND2X1 U7053 ( .A(n13834), .B(n13336), .Y(n13827) );
  INVX1 U7054 ( .A(n13827), .Y(n10499) );
  INVX1 U7055 ( .A(n10502), .Y(n10500) );
  INVX1 U7056 ( .A(n10500), .Y(n10501) );
  AND2X1 U7057 ( .A(n13371), .B(n13372), .Y(n13822) );
  INVX1 U7058 ( .A(n13822), .Y(n10502) );
  INVX1 U7059 ( .A(n10505), .Y(n10503) );
  INVX1 U7060 ( .A(n10503), .Y(n10504) );
  BUFX2 U7061 ( .A(n11677), .Y(n10505) );
  INVX1 U7062 ( .A(n10508), .Y(n10506) );
  INVX1 U7063 ( .A(n10506), .Y(n10507) );
  BUFX2 U7064 ( .A(n11955), .Y(n10508) );
  INVX1 U7065 ( .A(n10511), .Y(n10509) );
  INVX1 U7066 ( .A(n10509), .Y(n10510) );
  AND2X1 U7067 ( .A(\add_x_129/n1 ), .B(
        \lamb/scale_ts2/genblk1[3].mult/added[4] ), .Y(n11721) );
  INVX1 U7068 ( .A(n11721), .Y(n10511) );
  INVX1 U7069 ( .A(n10514), .Y(n10512) );
  INVX1 U7070 ( .A(n10512), .Y(n10513) );
  AND2X1 U7071 ( .A(\add_x_145/n1 ), .B(
        \lamb/scale_ts1/genblk1[0].mult/added[4] ), .Y(n12740) );
  INVX1 U7072 ( .A(n12740), .Y(n10514) );
  INVX1 U7073 ( .A(n10517), .Y(n10515) );
  INVX1 U7074 ( .A(n10515), .Y(n10516) );
  AND2X2 U7075 ( .A(n12391), .B(n12290), .Y(n12407) );
  INVX1 U7076 ( .A(n12407), .Y(n10517) );
  INVX1 U7077 ( .A(n10520), .Y(n10518) );
  INVX1 U7078 ( .A(n10518), .Y(n10519) );
  BUFX2 U7079 ( .A(n12243), .Y(n10520) );
  INVX1 U7080 ( .A(n10523), .Y(n10521) );
  INVX1 U7081 ( .A(n10521), .Y(n10522) );
  AND2X1 U7082 ( .A(\lamb/scale_ts3/genblk1[3].mult/added[1] ), .B(
        \lamb/scale_ts3/genblk1[3].mult/added[2] ), .Y(n12579) );
  INVX1 U7083 ( .A(n12579), .Y(n10523) );
  INVX1 U7084 ( .A(n10526), .Y(n10524) );
  INVX1 U7085 ( .A(n10524), .Y(n10525) );
  BUFX2 U7086 ( .A(n13564), .Y(n10526) );
  INVX1 U7087 ( .A(n10529), .Y(n10527) );
  INVX1 U7088 ( .A(n10527), .Y(n10528) );
  AND2X1 U7089 ( .A(n13225), .B(n13231), .Y(n12761) );
  INVX1 U7090 ( .A(n12761), .Y(n10529) );
  INVX1 U7091 ( .A(n10532), .Y(n10530) );
  INVX1 U7092 ( .A(n10530), .Y(n10531) );
  BUFX2 U7093 ( .A(n13566), .Y(n10532) );
  INVX1 U7094 ( .A(n10535), .Y(n10533) );
  INVX1 U7095 ( .A(n10533), .Y(n10534) );
  AND2X2 U7096 ( .A(n13424), .B(n13411), .Y(n13444) );
  INVX1 U7097 ( .A(n13444), .Y(n10535) );
  INVX1 U7098 ( .A(n10538), .Y(n10536) );
  INVX1 U7099 ( .A(n10536), .Y(n10537) );
  BUFX2 U7100 ( .A(n12543), .Y(n10538) );
  INVX1 U7101 ( .A(n10541), .Y(n10539) );
  INVX1 U7102 ( .A(n10539), .Y(n10540) );
  BUFX2 U7103 ( .A(n13533), .Y(n10541) );
  INVX1 U7104 ( .A(n10544), .Y(n10542) );
  INVX1 U7105 ( .A(n10542), .Y(n10543) );
  OR2X1 U7106 ( .A(n10678), .B(n10743), .Y(n13030) );
  INVX1 U7107 ( .A(n13030), .Y(n10544) );
  INVX1 U7108 ( .A(n10547), .Y(n10545) );
  INVX1 U7109 ( .A(n10545), .Y(n10546) );
  AND2X1 U7110 ( .A(n10793), .B(n12935), .Y(n12806) );
  INVX1 U7111 ( .A(n12806), .Y(n10547) );
  INVX1 U7112 ( .A(n10550), .Y(n10548) );
  INVX1 U7113 ( .A(n10548), .Y(n10549) );
  AND2X1 U7114 ( .A(n12690), .B(n13868), .Y(n13872) );
  INVX1 U7115 ( .A(n13872), .Y(n10550) );
  INVX1 U7116 ( .A(n10553), .Y(n10551) );
  INVX1 U7117 ( .A(n10551), .Y(n10552) );
  BUFX2 U7118 ( .A(n11452), .Y(n10553) );
  INVX1 U7119 ( .A(n10556), .Y(n10554) );
  INVX1 U7120 ( .A(n10554), .Y(n10555) );
  BUFX2 U7121 ( .A(n11846), .Y(n10556) );
  INVX1 U7122 ( .A(n10559), .Y(n10557) );
  INVX1 U7123 ( .A(n10557), .Y(n10558) );
  BUFX2 U7124 ( .A(n12499), .Y(n10559) );
  INVX1 U7125 ( .A(n10562), .Y(n10560) );
  INVX1 U7126 ( .A(n10560), .Y(n10561) );
  BUFX2 U7127 ( .A(n12520), .Y(n10562) );
  INVX1 U7128 ( .A(n10565), .Y(n10563) );
  INVX1 U7129 ( .A(n10563), .Y(n10564) );
  AND2X1 U7130 ( .A(n13903), .B(n12795), .Y(n12844) );
  INVX1 U7131 ( .A(n12844), .Y(n10565) );
  INVX1 U7132 ( .A(n10568), .Y(n10566) );
  INVX1 U7133 ( .A(n10566), .Y(n10567) );
  BUFX2 U7134 ( .A(n12979), .Y(n10568) );
  INVX1 U7135 ( .A(n10571), .Y(n10569) );
  INVX1 U7136 ( .A(n10569), .Y(n10570) );
  AND2X1 U7137 ( .A(n13489), .B(n12795), .Y(n12944) );
  INVX1 U7138 ( .A(n12944), .Y(n10571) );
  INVX1 U7139 ( .A(n10574), .Y(n10572) );
  INVX1 U7140 ( .A(n10572), .Y(n10573) );
  AND2X1 U7141 ( .A(n12431), .B(n13586), .Y(n13484) );
  INVX1 U7142 ( .A(n13484), .Y(n10574) );
  INVX1 U7143 ( .A(n10577), .Y(n10575) );
  INVX1 U7144 ( .A(n10575), .Y(n10576) );
  AND2X1 U7145 ( .A(n13903), .B(n10984), .Y(n13006) );
  INVX1 U7146 ( .A(n13006), .Y(n10577) );
  INVX1 U7147 ( .A(n10580), .Y(n10578) );
  INVX1 U7148 ( .A(n10578), .Y(n10579) );
  AND2X2 U7149 ( .A(n10828), .B(n12703), .Y(n13244) );
  INVX1 U7150 ( .A(n13244), .Y(n10580) );
  INVX1 U7151 ( .A(n10583), .Y(n10581) );
  INVX1 U7152 ( .A(n10581), .Y(n10582) );
  AND2X1 U7153 ( .A(n12152), .B(n12804), .Y(n12929) );
  INVX1 U7154 ( .A(n12929), .Y(n10583) );
  INVX1 U7155 ( .A(n10586), .Y(n10584) );
  INVX1 U7156 ( .A(n10584), .Y(n10585) );
  AND2X1 U7157 ( .A(n13439), .B(n13437), .Y(n13459) );
  INVX1 U7158 ( .A(n13459), .Y(n10586) );
  INVX1 U7159 ( .A(n10589), .Y(n10587) );
  INVX1 U7160 ( .A(n10587), .Y(n10588) );
  BUFX2 U7161 ( .A(n11990), .Y(n10589) );
  INVX1 U7162 ( .A(n10592), .Y(n10590) );
  INVX1 U7163 ( .A(n10590), .Y(n10591) );
  AND2X1 U7164 ( .A(n13840), .B(n13848), .Y(n12697) );
  INVX1 U7165 ( .A(n12697), .Y(n10592) );
  INVX1 U7166 ( .A(n10595), .Y(n10593) );
  INVX1 U7167 ( .A(n10593), .Y(n10594) );
  AND2X1 U7168 ( .A(n10849), .B(n13131), .Y(n13134) );
  INVX1 U7169 ( .A(n13134), .Y(n10595) );
  INVX1 U7170 ( .A(n10598), .Y(n10596) );
  INVX1 U7171 ( .A(n10596), .Y(n10597) );
  BUFX2 U7172 ( .A(n12595), .Y(n10598) );
  INVX1 U7173 ( .A(n10601), .Y(n10599) );
  INVX1 U7174 ( .A(n10599), .Y(n10600) );
  AND2X1 U7175 ( .A(n12724), .B(n12723), .Y(n13929) );
  INVX1 U7176 ( .A(n13929), .Y(n10601) );
  INVX1 U7177 ( .A(n10604), .Y(n10602) );
  INVX1 U7178 ( .A(n10602), .Y(n10603) );
  OR2X2 U7179 ( .A(n11651), .B(n11650), .Y(n11689) );
  INVX1 U7180 ( .A(n11689), .Y(n10604) );
  INVX1 U7181 ( .A(n10607), .Y(n10605) );
  INVX1 U7182 ( .A(n10605), .Y(n10606) );
  AND2X1 U7183 ( .A(n13085), .B(n12696), .Y(n12684) );
  INVX1 U7184 ( .A(n12684), .Y(n10607) );
  INVX1 U7185 ( .A(n10610), .Y(n10608) );
  INVX1 U7186 ( .A(n10608), .Y(n10609) );
  AND2X1 U7187 ( .A(n12787), .B(n11192), .Y(n13585) );
  INVX1 U7188 ( .A(n13585), .Y(n10610) );
  INVX1 U7189 ( .A(n10613), .Y(n10611) );
  INVX1 U7190 ( .A(n10611), .Y(n10612) );
  AND2X2 U7191 ( .A(n13752), .B(n12837), .Y(n12841) );
  INVX1 U7192 ( .A(n12841), .Y(n10613) );
  INVX1 U7193 ( .A(n10616), .Y(n10614) );
  INVX1 U7194 ( .A(n10614), .Y(n10615) );
  BUFX2 U7195 ( .A(n13508), .Y(n10616) );
  INVX1 U7196 ( .A(n10619), .Y(n10617) );
  INVX1 U7197 ( .A(n10617), .Y(n10618) );
  BUFX2 U7198 ( .A(n12301), .Y(n10619) );
  INVX1 U7199 ( .A(n10622), .Y(n10620) );
  INVX1 U7200 ( .A(n10620), .Y(n10621) );
  AND2X2 U7201 ( .A(n11476), .B(n11475), .Y(n11492) );
  INVX1 U7202 ( .A(n11492), .Y(n10622) );
  INVX1 U7203 ( .A(n10625), .Y(n10623) );
  INVX1 U7204 ( .A(n10623), .Y(n10624) );
  BUFX2 U7205 ( .A(n13543), .Y(n10625) );
  OR2X1 U7206 ( .A(n13371), .B(n11127), .Y(n13376) );
  OR2X1 U7207 ( .A(n10703), .B(n10800), .Y(n13943) );
  AND2X1 U7208 ( .A(n11558), .B(n10997), .Y(n11619) );
  OR2X1 U7209 ( .A(n11003), .B(n13917), .Y(n13217) );
  AND2X1 U7210 ( .A(n10734), .B(n11411), .Y(n11416) );
  XOR2X1 U7211 ( .A(n11010), .B(n10971), .Y(n13326) );
  OR2X1 U7212 ( .A(n12353), .B(n10917), .Y(n12355) );
  AND2X1 U7213 ( .A(n11327), .B(n11173), .Y(n11308) );
  OR2X1 U7214 ( .A(n10828), .B(n11169), .Y(n13249) );
  AND2X1 U7215 ( .A(n10994), .B(n11403), .Y(n11407) );
  OR2X1 U7216 ( .A(n11760), .B(n10629), .Y(n11548) );
  AND2X1 U7217 ( .A(n13151), .B(n10995), .Y(n13169) );
  OR2X1 U7218 ( .A(n12288), .B(n10634), .Y(n12391) );
  AND2X1 U7219 ( .A(n10634), .B(n12288), .Y(n12387) );
  OR2X1 U7220 ( .A(n11519), .B(n11048), .Y(n11523) );
  AND2X1 U7221 ( .A(n11195), .B(n10742), .Y(n12941) );
  AND2X1 U7222 ( .A(n11832), .B(n10752), .Y(n11855) );
  AND2X1 U7223 ( .A(n10678), .B(n10743), .Y(n13034) );
  AND2X1 U7224 ( .A(n12433), .B(n10667), .Y(n12545) );
  AND2X1 U7225 ( .A(n11174), .B(n10900), .Y(n13845) );
  OR2X1 U7226 ( .A(n10785), .B(n13912), .Y(n10364) );
  AND2X1 U7227 ( .A(n13062), .B(n11095), .Y(n13055) );
  AND2X1 U7228 ( .A(n12898), .B(n11207), .Y(n12779) );
  AND2X1 U7229 ( .A(n11176), .B(n10989), .Y(n12976) );
  AND2X1 U7230 ( .A(n12984), .B(n11176), .Y(n12980) );
  OR2X1 U7231 ( .A(n11203), .B(n12829), .Y(n12810) );
  AND2X1 U7232 ( .A(n12853), .B(n10793), .Y(n13588) );
  OR2X1 U7233 ( .A(n11203), .B(n12855), .Y(n12856) );
  OR2X1 U7234 ( .A(n10727), .B(n13891), .Y(n12970) );
  OR2X1 U7235 ( .A(n11140), .B(n10782), .Y(n13540) );
  AND2X1 U7236 ( .A(n12905), .B(n12867), .Y(n12868) );
  OR2X1 U7237 ( .A(n11192), .B(n12432), .Y(n12862) );
  AND2X1 U7238 ( .A(n10725), .B(n12975), .Y(n12988) );
  AND2X1 U7239 ( .A(n10680), .B(n10742), .Y(n12922) );
  OR2X1 U7240 ( .A(n11327), .B(n10669), .Y(n11310) );
  OR2X1 U7241 ( .A(n11788), .B(n10641), .Y(n11789) );
  AND2X1 U7242 ( .A(n13258), .B(n10630), .Y(n13218) );
  AND2X1 U7243 ( .A(n10629), .B(n11760), .Y(n11761) );
  AND2X1 U7244 ( .A(n13342), .B(n12292), .Y(n13873) );
  INVX1 U7245 ( .A(n13873), .Y(n10626) );
  AND2X1 U7246 ( .A(n10851), .B(n11714), .Y(n13258) );
  INVX1 U7247 ( .A(n13258), .Y(n10627) );
  OR2X1 U7248 ( .A(n12448), .B(\lamb/scale_ds2/genblk1[2].mult/added[3] ), .Y(
        n12481) );
  INVX1 U7249 ( .A(n12481), .Y(n10628) );
  OR2X1 U7250 ( .A(\lamb/scale_ds2/genblk1[3].mult/added[4] ), .B(
        \add_x_133/n1 ), .Y(n11550) );
  INVX1 U7251 ( .A(n11550), .Y(n10629) );
  AND2X1 U7252 ( .A(n12673), .B(n12672), .Y(n13381) );
  INVX1 U7253 ( .A(n13381), .Y(n10630) );
  BUFX2 U7254 ( .A(n12360), .Y(n10631) );
  OR2X1 U7255 ( .A(n13702), .B(n10729), .Y(n13772) );
  INVX1 U7256 ( .A(n13772), .Y(n10632) );
  AND2X1 U7257 ( .A(n13567), .B(n13556), .Y(n13643) );
  INVX1 U7258 ( .A(n13643), .Y(n10633) );
  OR2X1 U7259 ( .A(\add_x_117/n1 ), .B(
        \lamb/scale_ts3/genblk1[2].mult/added[4] ), .Y(n12375) );
  INVX1 U7260 ( .A(n12375), .Y(n10634) );
  AND2X1 U7261 ( .A(n12695), .B(n12682), .Y(n11713) );
  INVX1 U7262 ( .A(n11713), .Y(n10635) );
  OR2X1 U7263 ( .A(n10728), .B(n10730), .Y(n13773) );
  INVX1 U7264 ( .A(n13773), .Y(n10636) );
  BUFX2 U7265 ( .A(n11754), .Y(n10637) );
  OR2X1 U7266 ( .A(n13650), .B(n13613), .Y(n13759) );
  INVX1 U7267 ( .A(n13759), .Y(n10638) );
  OR2X1 U7268 ( .A(n13635), .B(n13650), .Y(n13762) );
  INVX1 U7269 ( .A(n13762), .Y(n10639) );
  BUFX2 U7270 ( .A(n13469), .Y(n10640) );
  AND2X1 U7271 ( .A(\lamb/scale_bs3/genblk1[0].mult/added[4] ), .B(
        \add_x_125/n1 ), .Y(n11787) );
  INVX1 U7272 ( .A(n11787), .Y(n10641) );
  AND2X1 U7273 ( .A(\lamb/scale_ts0/genblk1[1].mult/added[2] ), .B(
        \lamb/scale_ts0/genblk1[1].mult/added[1] ), .Y(n11620) );
  INVX1 U7274 ( .A(n11620), .Y(n10642) );
  AND2X1 U7275 ( .A(\lamb/scale_ls2/genblk1[1].mult/added[3] ), .B(n11830), 
        .Y(n11835) );
  INVX1 U7276 ( .A(n11835), .Y(n10643) );
  BUFX2 U7277 ( .A(n13405), .Y(n10644) );
  AND2X1 U7278 ( .A(\lamb/scale_ts2/genblk1[2].mult/added[1] ), .B(
        \lamb/scale_ts2/genblk1[2].mult/added[2] ), .Y(n12483) );
  INVX1 U7279 ( .A(n12483), .Y(n10645) );
  AND2X1 U7280 ( .A(n12752), .B(n11003), .Y(n13913) );
  INVX1 U7281 ( .A(n13913), .Y(n10646) );
  BUFX2 U7282 ( .A(n13569), .Y(n10647) );
  BUFX2 U7283 ( .A(n13560), .Y(n10648) );
  AND2X1 U7284 ( .A(\forney/m1/added [4]), .B(\add_x_20/n1 ), .Y(n13496) );
  INVX1 U7285 ( .A(n13496), .Y(n10649) );
  AND2X1 U7286 ( .A(n13077), .B(n13072), .Y(n13073) );
  INVX1 U7287 ( .A(n13073), .Y(n10650) );
  AND2X1 U7288 ( .A(n13053), .B(n13061), .Y(n13054) );
  INVX1 U7289 ( .A(n13054), .Y(n10651) );
  AND2X1 U7290 ( .A(n12222), .B(n12254), .Y(n12274) );
  INVX1 U7291 ( .A(n12274), .Y(n10652) );
  AND2X1 U7292 ( .A(\lamb/scale_ts1/genblk1[1].mult/added[3] ), .B(n12296), 
        .Y(n12351) );
  INVX1 U7293 ( .A(n12351), .Y(n10653) );
  BUFX2 U7294 ( .A(n11899), .Y(n10654) );
  AND2X1 U7295 ( .A(n13547), .B(n13535), .Y(n13529) );
  INVX1 U7296 ( .A(n13529), .Y(n10655) );
  BUFX2 U7297 ( .A(n11378), .Y(n10656) );
  AND2X1 U7298 ( .A(n11075), .B(n10808), .Y(n13286) );
  INVX1 U7299 ( .A(n13286), .Y(n10657) );
  INVX1 U7300 ( .A(n13041), .Y(n10658) );
  AND2X1 U7301 ( .A(n11163), .B(n10612), .Y(n13005) );
  INVX1 U7302 ( .A(n13005), .Y(n10659) );
  AND2X1 U7303 ( .A(n11159), .B(n11475), .Y(n11493) );
  INVX1 U7304 ( .A(n11493), .Y(n10660) );
  AND2X1 U7305 ( .A(\forney/pe0/mult0/added [3]), .B(n12572), .Y(n12531) );
  INVX1 U7306 ( .A(n12531), .Y(n10661) );
  OR2X1 U7307 ( .A(n13424), .B(n13443), .Y(n13454) );
  INVX1 U7308 ( .A(n13454), .Y(n10662) );
  AND2X1 U7309 ( .A(n12206), .B(n11184), .Y(n12204) );
  INVX1 U7310 ( .A(n12204), .Y(n10663) );
  AND2X1 U7311 ( .A(n13590), .B(n12848), .Y(n13593) );
  INVX1 U7312 ( .A(n13593), .Y(n10664) );
  AND2X1 U7313 ( .A(n12827), .B(n12935), .Y(n13750) );
  INVX1 U7314 ( .A(n13750), .Y(n10665) );
  OR2X1 U7315 ( .A(n11419), .B(\lamb/scale_ts1/genblk1[3].mult/added[3] ), .Y(
        n11417) );
  INVX1 U7316 ( .A(n11417), .Y(n10666) );
  AND2X1 U7317 ( .A(\lamb/scale_ds3/genblk1[3].mult/added[3] ), .B(n12547), 
        .Y(n12541) );
  INVX1 U7318 ( .A(n12541), .Y(n10667) );
  OR2X1 U7319 ( .A(n11304), .B(\add_x_146/n1 ), .Y(n11431) );
  INVX1 U7320 ( .A(n11431), .Y(n10668) );
  AND2X1 U7321 ( .A(\lamb/scale_ts0/genblk1[2].mult/added[4] ), .B(
        \add_x_152/n1 ), .Y(n11326) );
  INVX1 U7322 ( .A(n11326), .Y(n10669) );
  BUFX2 U7323 ( .A(n11525), .Y(n10670) );
  AND2X1 U7324 ( .A(n10609), .B(n11195), .Y(n12962) );
  INVX1 U7325 ( .A(n12962), .Y(n10671) );
  AND2X1 U7326 ( .A(\lamb/scale_ts1/genblk1[3].mult/added[3] ), .B(n11404), 
        .Y(n11406) );
  INVX1 U7327 ( .A(n11406), .Y(n10672) );
  BUFX2 U7328 ( .A(n13107), .Y(n10673) );
  AND2X1 U7329 ( .A(n10606), .B(n11174), .Y(n13314) );
  INVX1 U7330 ( .A(n13314), .Y(n10674) );
  BUFX2 U7331 ( .A(n11989), .Y(n10675) );
  BUFX2 U7332 ( .A(n12514), .Y(n10676) );
  AND2X1 U7333 ( .A(n13147), .B(n13138), .Y(n11995) );
  INVX1 U7334 ( .A(n11995), .Y(n10677) );
  BUFX2 U7335 ( .A(n12624), .Y(n10678) );
  BUFX2 U7336 ( .A(n11779), .Y(n10679) );
  AND2X1 U7337 ( .A(n13586), .B(n13590), .Y(n12827) );
  INVX1 U7338 ( .A(n12827), .Y(n10680) );
  BUFX2 U7339 ( .A(n13288), .Y(n10681) );
  AND2X1 U7340 ( .A(\add_x_117/n1 ), .B(
        \lamb/scale_ts3/genblk1[2].mult/added[4] ), .Y(n12289) );
  INVX1 U7341 ( .A(n12289), .Y(n10682) );
  INVX1 U7342 ( .A(n10683), .Y(n12905) );
  INVX1 U7343 ( .A(n12864), .Y(n10684) );
  INVX1 U7344 ( .A(n12865), .Y(n10685) );
  INVX1 U7345 ( .A(n12866), .Y(n10686) );
  NOR2X1 U7346 ( .A(n10686), .B(n10687), .Y(n10683) );
  NOR2X1 U7347 ( .A(n10684), .B(n10685), .Y(n10688) );
  INVX1 U7348 ( .A(n10688), .Y(n10687) );
  AND2X1 U7349 ( .A(n11712), .B(n11474), .Y(n12678) );
  INVX1 U7350 ( .A(n12678), .Y(n10689) );
  BUFX2 U7351 ( .A(n13045), .Y(n10690) );
  BUFX2 U7352 ( .A(n13485), .Y(n10691) );
  BUFX2 U7353 ( .A(n11248), .Y(n10692) );
  BUFX2 U7354 ( .A(n11290), .Y(n10693) );
  BUFX2 U7355 ( .A(n11352), .Y(n10694) );
  BUFX2 U7356 ( .A(n11396), .Y(n10695) );
  BUFX2 U7357 ( .A(n12647), .Y(n10696) );
  BUFX2 U7358 ( .A(n13472), .Y(n10697) );
  OR2X1 U7359 ( .A(n10753), .B(n13602), .Y(n13600) );
  INVX1 U7360 ( .A(n13600), .Y(n10698) );
  AND2X1 U7361 ( .A(n12431), .B(n12833), .Y(n13483) );
  INVX1 U7362 ( .A(n13483), .Y(n10699) );
  BUFX2 U7363 ( .A(n11499), .Y(n10700) );
  BUFX2 U7364 ( .A(n10377), .Y(n10701) );
  AND2X1 U7365 ( .A(\lamb/scale_ts0/genblk1[0].mult/added[1] ), .B(
        \lamb/scale_ts0/genblk1[0].mult/added[2] ), .Y(n12201) );
  INVX1 U7366 ( .A(n12201), .Y(n10702) );
  BUFX2 U7367 ( .A(n13187), .Y(n10703) );
  OR2X1 U7368 ( .A(n10730), .B(n11170), .Y(n13777) );
  INVX1 U7369 ( .A(n13777), .Y(n10704) );
  OR2X1 U7370 ( .A(n10730), .B(n10740), .Y(n13781) );
  INVX1 U7371 ( .A(n13781), .Y(n10705) );
  OR2X1 U7372 ( .A(n10730), .B(n13712), .Y(n13785) );
  INVX1 U7373 ( .A(n13785), .Y(n10706) );
  OR2X1 U7374 ( .A(n10728), .B(n10741), .Y(n13805) );
  INVX1 U7375 ( .A(n13805), .Y(n10707) );
  OR2X1 U7376 ( .A(n11170), .B(n10741), .Y(n13809) );
  INVX1 U7377 ( .A(n13809), .Y(n10708) );
  OR2X1 U7378 ( .A(n10740), .B(n10741), .Y(n13813) );
  INVX1 U7379 ( .A(n13813), .Y(n10709) );
  OR2X1 U7380 ( .A(n13712), .B(n10741), .Y(n13819) );
  INVX1 U7381 ( .A(n13819), .Y(n10710) );
  OR2X1 U7382 ( .A(n10729), .B(n13759), .Y(n13776) );
  INVX1 U7383 ( .A(n13776), .Y(n10711) );
  OR2X1 U7384 ( .A(n10729), .B(n13762), .Y(n13780) );
  INVX1 U7385 ( .A(n13780), .Y(n10712) );
  OR2X1 U7386 ( .A(n10729), .B(n13713), .Y(n13784) );
  INVX1 U7387 ( .A(n13784), .Y(n10713) );
  OR2X1 U7388 ( .A(n13702), .B(n11171), .Y(n13788) );
  INVX1 U7389 ( .A(n13788), .Y(n10714) );
  OR2X1 U7390 ( .A(n13759), .B(n11171), .Y(n13792) );
  INVX1 U7391 ( .A(n13792), .Y(n10715) );
  OR2X1 U7392 ( .A(n13762), .B(n11171), .Y(n13796) );
  INVX1 U7393 ( .A(n13796), .Y(n10716) );
  OR2X1 U7394 ( .A(n13713), .B(n11171), .Y(n13800) );
  INVX1 U7395 ( .A(n13800), .Y(n10717) );
  INVX1 U7396 ( .A(n10718), .Y(n13443) );
  INVX1 U7397 ( .A(n13394), .Y(n10719) );
  INVX1 U7398 ( .A(n13421), .Y(n10720) );
  NOR2X1 U7399 ( .A(n10720), .B(n10721), .Y(n10718) );
  NOR2X1 U7400 ( .A(n13393), .B(n10719), .Y(n10722) );
  INVX1 U7401 ( .A(n10722), .Y(n10721) );
  AND2X1 U7402 ( .A(n12682), .B(n13385), .Y(n11622) );
  INVX1 U7403 ( .A(n11622), .Y(n10723) );
  OR2X1 U7404 ( .A(n12225), .B(n12224), .Y(n13070) );
  INVX1 U7405 ( .A(n13070), .Y(n10724) );
  BUFX2 U7406 ( .A(n12977), .Y(n10725) );
  BUFX2 U7407 ( .A(n13175), .Y(n10726) );
  AND2X1 U7408 ( .A(n13488), .B(n12803), .Y(n13489) );
  INVX1 U7409 ( .A(n13489), .Y(n10727) );
  AND2X1 U7410 ( .A(n13662), .B(n13573), .Y(n13689) );
  INVX1 U7411 ( .A(n13689), .Y(n10728) );
  AND2X1 U7412 ( .A(n13574), .B(n13753), .Y(n13654) );
  INVX1 U7413 ( .A(n13654), .Y(n10729) );
  AND2X1 U7414 ( .A(n13748), .B(n13675), .Y(n13664) );
  INVX1 U7415 ( .A(n13664), .Y(n10730) );
  OR2X1 U7416 ( .A(\add_x_124/n1 ), .B(
        \lamb/scale_bs3/genblk1[1].mult/added[4] ), .Y(n11968) );
  INVX1 U7417 ( .A(n11968), .Y(n10731) );
  BUFX2 U7418 ( .A(n13869), .Y(n10732) );
  BUFX2 U7419 ( .A(n13039), .Y(n10733) );
  AND2X1 U7420 ( .A(\lamb/scale_ts1/genblk1[3].mult/added[3] ), .B(n11419), 
        .Y(n11412) );
  INVX1 U7421 ( .A(n11412), .Y(n10734) );
  INVX1 U7422 ( .A(n10735), .Y(n13712) );
  INVX1 U7423 ( .A(n13662), .Y(n10736) );
  INVX1 U7424 ( .A(n13663), .Y(n10737) );
  NOR2X1 U7425 ( .A(n10737), .B(n10738), .Y(n10735) );
  NOR2X1 U7426 ( .A(n13661), .B(n10736), .Y(n10739) );
  INVX1 U7427 ( .A(n10739), .Y(n10738) );
  AND2X1 U7428 ( .A(n13494), .B(n13493), .Y(n13662) );
  AND2X1 U7429 ( .A(n13662), .B(n13644), .Y(n13709) );
  INVX1 U7430 ( .A(n13709), .Y(n10740) );
  AND2X1 U7431 ( .A(n11175), .B(n13748), .Y(n13685) );
  INVX1 U7432 ( .A(n13685), .Y(n10741) );
  AND2X1 U7433 ( .A(n12826), .B(n10798), .Y(n13690) );
  INVX1 U7434 ( .A(n13690), .Y(n10742) );
  BUFX2 U7435 ( .A(n13025), .Y(n10743) );
  INVX1 U7436 ( .A(n10744), .Y(n13925) );
  INVX1 U7437 ( .A(n13927), .Y(n10745) );
  INVX1 U7438 ( .A(n12213), .Y(n10746) );
  NOR2X1 U7439 ( .A(n10746), .B(n10747), .Y(n10744) );
  NOR2X1 U7440 ( .A(n10745), .B(n12212), .Y(n10748) );
  INVX1 U7441 ( .A(n10748), .Y(n10747) );
  AND2X1 U7442 ( .A(n12760), .B(n12685), .Y(n12762) );
  INVX1 U7443 ( .A(n12762), .Y(n10749) );
  OR2X1 U7444 ( .A(n12627), .B(n13015), .Y(n13021) );
  INVX1 U7445 ( .A(n13021), .Y(n10750) );
  AND2X1 U7446 ( .A(\lamb/scale_ts1/genblk1[0].mult/added[1] ), .B(
        \lamb/scale_ts1/genblk1[0].mult/added[2] ), .Y(n12753) );
  INVX1 U7447 ( .A(n12753), .Y(n10751) );
  AND2X1 U7448 ( .A(\lamb/scale_ls2/genblk1[1].mult/added[3] ), .B(n11823), 
        .Y(n11837) );
  INVX1 U7449 ( .A(n11837), .Y(n10752) );
  AND2X1 U7450 ( .A(n12823), .B(n12930), .Y(n13744) );
  INVX1 U7451 ( .A(n13744), .Y(n10753) );
  AND2X1 U7452 ( .A(\lamb/scale_ds1/genblk1[1].mult/added[2] ), .B(
        \lamb/scale_ds1/genblk1[1].mult/added[1] ), .Y(n12339) );
  INVX1 U7453 ( .A(n12339), .Y(n10754) );
  BUFX2 U7454 ( .A(n12648), .Y(n10755) );
  BUFX2 U7455 ( .A(\lamb/scale_ds2/genblk1[3].mult/logA[1] ), .Y(n10756) );
  BUFX2 U7456 ( .A(n10361), .Y(n10757) );
  BUFX2 U7457 ( .A(\lamb/scale_ds3/genblk1[3].mult/logA[2] ), .Y(n10758) );
  BUFX2 U7458 ( .A(\forney/m0/logA [0]), .Y(n10759) );
  BUFX2 U7459 ( .A(\lamb/scale_ds3/genblk1[2].mult/logA[1] ), .Y(n10760) );
  BUFX2 U7460 ( .A(\lamb/scale_ds3/genblk1[2].mult/logA[2] ), .Y(n10761) );
  BUFX2 U7461 ( .A(\lamb/scale_ls3/genblk1[2].mult/logA[0] ), .Y(n10762) );
  OR2X1 U7462 ( .A(n12629), .B(n10750), .Y(\forney/pe0/mult0/logA [0]) );
  BUFX2 U7463 ( .A(\lamb/scale_ls3/genblk1[1].mult/logA[2] ), .Y(n10763) );
  BUFX2 U7464 ( .A(\lamb/scale_ls3/genblk1[0].mult/logA[1] ), .Y(n10764) );
  BUFX2 U7465 ( .A(\lamb/scale_ts2/genblk1[1].mult/logA[1] ), .Y(n10765) );
  BUFX2 U7466 ( .A(\lamb/scale_ds2/genblk1[2].mult/logA[1] ), .Y(n10766) );
  BUFX2 U7467 ( .A(\lamb/scale_ds2/genblk1[1].mult/logA[1] ), .Y(n10767) );
  BUFX2 U7468 ( .A(\lamb/scale_bs2/genblk1[0].mult/logA[2] ), .Y(n10768) );
  BUFX2 U7469 ( .A(\lamb/scale_ts1/genblk1[2].mult/logA[1] ), .Y(n10769) );
  BUFX2 U7470 ( .A(\lamb/scale_ts1/genblk1[2].mult/logA[2] ), .Y(n10770) );
  BUFX2 U7471 ( .A(\lamb/scale_ts1/genblk1[1].mult/logA[2] ), .Y(n10771) );
  BUFX2 U7472 ( .A(\lamb/scale_ds1/genblk1[3].mult/logA[1] ), .Y(n10772) );
  BUFX2 U7473 ( .A(\lamb/scale_ds1/genblk1[2].mult/logA[2] ), .Y(n10773) );
  BUFX2 U7474 ( .A(\lamb/scale_ts0/genblk1[1].mult/logA[1] ), .Y(n10774) );
  BUFX2 U7475 ( .A(n10373), .Y(n10775) );
  BUFX2 U7476 ( .A(n10369), .Y(n10776) );
  BUFX2 U7477 ( .A(n10366), .Y(n10777) );
  INVX1 U7478 ( .A(\lamb/scale_bs3/genblk1[1].mult/logA[1] ), .Y(n10778) );
  OR2X1 U7479 ( .A(n13844), .B(n12764), .Y(
        \lamb/scale_bs3/genblk1[1].mult/logA[1] ) );
  INVX1 U7480 ( .A(\lamb/scale_ls3/genblk1[0].mult/logA[0] ), .Y(n10779) );
  AND2X1 U7481 ( .A(n12770), .B(n11177), .Y(
        \lamb/scale_ls3/genblk1[0].mult/logA[0] ) );
  INVX1 U7482 ( .A(\lamb/scale_ls3/genblk1[2].mult/logA[1] ), .Y(n10780) );
  OR2X1 U7483 ( .A(n11136), .B(n13111), .Y(
        \lamb/scale_ls3/genblk1[2].mult/logA[1] ) );
  INVX1 U7484 ( .A(\lamb/scale_ts2/genblk1[3].mult/logA[1] ), .Y(n10781) );
  OR2X1 U7485 ( .A(n11023), .B(n13156), .Y(
        \lamb/scale_ts2/genblk1[3].mult/logA[1] ) );
  INVX1 U7486 ( .A(n13553), .Y(n10782) );
  OR2X1 U7487 ( .A(n10624), .B(n13542), .Y(n13553) );
  INVX1 U7488 ( .A(n11526), .Y(n10783) );
  AND2X1 U7489 ( .A(n11478), .B(\lamb/scale_ls2/genblk1[0].mult/added[3] ), 
        .Y(n11526) );
  BUFX2 U7490 ( .A(n12754), .Y(n10784) );
  INVX1 U7491 ( .A(n10365), .Y(n10785) );
  AND2X1 U7492 ( .A(n13911), .B(n13910), .Y(n10365) );
  BUFX2 U7493 ( .A(\lamb/scale_ts0/genblk1[0].mult/logA[2] ), .Y(n10786) );
  INVX1 U7494 ( .A(\lamb/scale_ts0/genblk1[0].mult/logA[1] ), .Y(n10787) );
  OR2X1 U7495 ( .A(n12673), .B(n12672), .Y(
        \lamb/scale_ts0/genblk1[0].mult/logA[1] ) );
  BUFX2 U7496 ( .A(\forney/m1/logB [1]), .Y(n10788) );
  BUFX2 U7497 ( .A(\forney/pe1/mult0/logB [1]), .Y(n10789) );
  BUFX2 U7498 ( .A(\forney/pe0/mult0/logB [1]), .Y(n10790) );
  BUFX2 U7499 ( .A(\forney/m1/logA [1]), .Y(n10791) );
  BUFX2 U7500 ( .A(n10378), .Y(n10792) );
  INVX1 U7501 ( .A(n12787), .Y(n10793) );
  AND2X1 U7502 ( .A(n12033), .B(n12032), .Y(n12787) );
  INVX1 U7503 ( .A(n10795), .Y(n10794) );
  BUFX2 U7504 ( .A(n13284), .Y(n10795) );
  INVX1 U7505 ( .A(n10797), .Y(n10796) );
  BUFX2 U7506 ( .A(n13289), .Y(n10797) );
  INVX1 U7507 ( .A(n13590), .Y(n10798) );
  AND2X1 U7508 ( .A(n12431), .B(n12771), .Y(n13590) );
  INVX1 U7509 ( .A(n11857), .Y(n10799) );
  AND2X1 U7510 ( .A(n12682), .B(n11024), .Y(n11857) );
  BUFX2 U7511 ( .A(n13186), .Y(n10800) );
  NOR2X1 U7512 ( .A(n10801), .B(n10802), .Y(n13186) );
  NOR2X1 U7513 ( .A(n11075), .B(n10809), .Y(n10801) );
  INVX1 U7514 ( .A(n13359), .Y(n10803) );
  NOR2X1 U7515 ( .A(n13235), .B(n10803), .Y(n10802) );
  INVX1 U7516 ( .A(n10805), .Y(n10804) );
  BUFX2 U7517 ( .A(n13188), .Y(n10805) );
  NOR2X1 U7518 ( .A(n10806), .B(n10807), .Y(n13188) );
  INVX1 U7519 ( .A(n10681), .Y(n10808) );
  INVX1 U7520 ( .A(n13235), .Y(n10809) );
  NOR2X1 U7521 ( .A(n10808), .B(n10809), .Y(n10806) );
  INVX1 U7522 ( .A(n10468), .Y(n10810) );
  NOR2X1 U7523 ( .A(n13235), .B(n10810), .Y(n10807) );
  INVX1 U7524 ( .A(n13630), .Y(n10811) );
  AND2X1 U7525 ( .A(n13605), .B(n13609), .Y(n13630) );
  INVX1 U7526 ( .A(n10813), .Y(n10812) );
  BUFX2 U7527 ( .A(n13028), .Y(n10813) );
  INVX1 U7528 ( .A(n10815), .Y(n10814) );
  BUFX2 U7529 ( .A(n11517), .Y(n10815) );
  INVX1 U7530 ( .A(n10817), .Y(n10816) );
  BUFX2 U7531 ( .A(n13178), .Y(n10817) );
  INVX1 U7532 ( .A(n13238), .Y(n10818) );
  AND2X1 U7533 ( .A(n13231), .B(n12696), .Y(n13238) );
  INVX1 U7534 ( .A(n10820), .Y(n10819) );
  BUFX2 U7535 ( .A(n13150), .Y(n10820) );
  INVX1 U7536 ( .A(n12083), .Y(n10821) );
  AND2X1 U7537 ( .A(n10585), .B(n13430), .Y(n12083) );
  INVX1 U7538 ( .A(n13081), .Y(n10822) );
  OR2X1 U7539 ( .A(n12282), .B(n12281), .Y(n13081) );
  INVX1 U7540 ( .A(n10824), .Y(n10823) );
  BUFX2 U7541 ( .A(n13132), .Y(n10824) );
  INVX1 U7542 ( .A(n11485), .Y(n10825) );
  OR2X1 U7543 ( .A(\add_x_138/n1 ), .B(
        \lamb/scale_bs2/genblk1[0].mult/added[4] ), .Y(n11485) );
  INVX1 U7544 ( .A(n13240), .Y(n10826) );
  AND2X1 U7545 ( .A(n13225), .B(n13224), .Y(n13240) );
  INVX1 U7546 ( .A(n10828), .Y(n10827) );
  BUFX2 U7547 ( .A(n13243), .Y(n10828) );
  INVX1 U7548 ( .A(n10830), .Y(n10829) );
  BUFX2 U7549 ( .A(n13046), .Y(n10830) );
  INVX1 U7550 ( .A(n10832), .Y(n10831) );
  BUFX2 U7551 ( .A(n13946), .Y(n10832) );
  INVX1 U7552 ( .A(n13752), .Y(n10833) );
  AND2X1 U7553 ( .A(n12964), .B(n11135), .Y(n13752) );
  BUFX2 U7554 ( .A(\lamb/scale_ls3/genblk1[0].mult/logB[3] ), .Y(n10834) );
  NAND2X1 U7555 ( .A(n10835), .B(n10836), .Y(
        \lamb/scale_ls3/genblk1[0].mult/logB[3] ) );
  INVX1 U7556 ( .A(n12702), .Y(n10837) );
  INVX1 U7557 ( .A(n13129), .Y(n10838) );
  NAND2X1 U7558 ( .A(n10837), .B(n10838), .Y(n10835) );
  NAND2X1 U7559 ( .A(n10837), .B(n10823), .Y(n10836) );
  INVX1 U7560 ( .A(n10840), .Y(n10839) );
  BUFX2 U7561 ( .A(n12058), .Y(n10840) );
  BUFX2 U7562 ( .A(\lamb/scale_ls2/genblk1[0].mult/logB[3] ), .Y(n10841) );
  BUFX2 U7563 ( .A(n12071), .Y(n10842) );
  BUFX2 U7564 ( .A(n12073), .Y(n10843) );
  BUFX2 U7565 ( .A(\lamb/scale_ls3/genblk1[0].mult/logB[1] ), .Y(n10844) );
  NOR2X1 U7566 ( .A(n10845), .B(n10846), .Y(
        \lamb/scale_ls3/genblk1[0].mult/logB[1] ) );
  INVX1 U7567 ( .A(n12709), .Y(n10847) );
  NOR2X1 U7568 ( .A(n10847), .B(n10823), .Y(n10845) );
  INVX1 U7569 ( .A(n12707), .Y(n10848) );
  INVX1 U7570 ( .A(n12708), .Y(n10849) );
  NOR2X1 U7571 ( .A(n10848), .B(n10849), .Y(n10846) );
  BUFX2 U7572 ( .A(\lamb/scale_ls2/genblk1[0].mult/logB[1] ), .Y(n10850) );
  INVX1 U7573 ( .A(n12682), .Y(n10851) );
  OR2X1 U7574 ( .A(n11394), .B(n10606), .Y(n12682) );
  INVX1 U7575 ( .A(n10852), .Y(n12913) );
  INVX1 U7576 ( .A(n12920), .Y(n10853) );
  INVX1 U7577 ( .A(n13492), .Y(n10854) );
  NOR2X1 U7578 ( .A(n10854), .B(n10855), .Y(n10852) );
  NOR2X1 U7579 ( .A(n13490), .B(n10853), .Y(n10856) );
  INVX1 U7580 ( .A(n10856), .Y(n10855) );
  INVX1 U7581 ( .A(n10857), .Y(n11642) );
  INVX1 U7582 ( .A(n10397), .Y(n10858) );
  INVX1 U7583 ( .A(n11641), .Y(n10859) );
  NOR2X1 U7584 ( .A(n10859), .B(n10860), .Y(n10857) );
  NOR2X1 U7585 ( .A(n10858), .B(\lamb/scale_ts1/genblk1[2].mult/added[3] ), 
        .Y(n10861) );
  INVX1 U7586 ( .A(n10861), .Y(n10860) );
  INVX1 U7587 ( .A(n10862), .Y(n13607) );
  INVX1 U7588 ( .A(n13631), .Y(n10863) );
  NOR2X1 U7589 ( .A(n13627), .B(n10864), .Y(n10862) );
  NOR2X1 U7590 ( .A(n10863), .B(n13630), .Y(n10865) );
  INVX1 U7591 ( .A(n10865), .Y(n10864) );
  BUFX2 U7592 ( .A(n12066), .Y(n10866) );
  BUFX2 U7593 ( .A(n12022), .Y(n10867) );
  BUFX2 U7594 ( .A(n12119), .Y(n10868) );
  BUFX2 U7595 ( .A(n12054), .Y(n10869) );
  BUFX2 U7596 ( .A(n12100), .Y(n10870) );
  XOR2X1 U7597 ( .A(n12110), .B(n12096), .Y(n12126) );
  BUFX2 U7598 ( .A(n12006), .Y(n10871) );
  AND2X1 U7599 ( .A(n10615), .B(n13507), .Y(n13501) );
  INVX1 U7600 ( .A(n13501), .Y(n10872) );
  AND2X1 U7601 ( .A(n12932), .B(n12819), .Y(n12820) );
  INVX1 U7602 ( .A(n12820), .Y(n10873) );
  BUFX2 U7603 ( .A(n13084), .Y(n10874) );
  INVX1 U7604 ( .A(n10875), .Y(n12453) );
  INVX1 U7605 ( .A(n12504), .Y(n10876) );
  INVX1 U7606 ( .A(\lamb/scale_ds2/genblk1[2].mult/added[2] ), .Y(n10877) );
  NOR2X1 U7607 ( .A(n10877), .B(n10878), .Y(n10875) );
  NOR2X1 U7608 ( .A(n10628), .B(n10876), .Y(n10879) );
  INVX1 U7609 ( .A(n10879), .Y(n10878) );
  BUFX2 U7610 ( .A(n12087), .Y(n10880) );
  INVX1 U7611 ( .A(n10881), .Y(n12902) );
  INVX1 U7612 ( .A(n12899), .Y(n10882) );
  INVX1 U7613 ( .A(n12900), .Y(n10883) );
  INVX1 U7614 ( .A(n12901), .Y(n10884) );
  NOR2X1 U7615 ( .A(n10884), .B(n10885), .Y(n10881) );
  NOR2X1 U7616 ( .A(n10882), .B(n10883), .Y(n10886) );
  INVX1 U7617 ( .A(n10886), .Y(n10885) );
  INVX1 U7618 ( .A(n10887), .Y(n11448) );
  INVX1 U7619 ( .A(n11446), .Y(n10888) );
  INVX1 U7620 ( .A(n11447), .Y(n10889) );
  NOR2X1 U7621 ( .A(n11442), .B(n10890), .Y(n10887) );
  NOR2X1 U7622 ( .A(n10888), .B(n10889), .Y(n10891) );
  INVX1 U7623 ( .A(n10891), .Y(n10890) );
  INVX1 U7624 ( .A(n10892), .Y(n12260) );
  INVX1 U7625 ( .A(n12257), .Y(n10893) );
  INVX1 U7626 ( .A(n12258), .Y(n10894) );
  INVX1 U7627 ( .A(n12259), .Y(n10895) );
  NOR2X1 U7628 ( .A(n10895), .B(n10896), .Y(n10892) );
  NOR2X1 U7629 ( .A(n10893), .B(n10894), .Y(n10897) );
  INVX1 U7630 ( .A(n10897), .Y(n10896) );
  AND2X1 U7631 ( .A(n11361), .B(n11360), .Y(n11362) );
  INVX1 U7632 ( .A(n11362), .Y(n10898) );
  BUFX2 U7633 ( .A(n13420), .Y(n10899) );
  AND2X1 U7634 ( .A(n13421), .B(n10899), .Y(n13450) );
  AND2X1 U7635 ( .A(n12696), .B(n12688), .Y(n12683) );
  INVX1 U7636 ( .A(n12683), .Y(n10900) );
  INVX1 U7637 ( .A(n10901), .Y(n11403) );
  INVX1 U7638 ( .A(\lamb/scale_ts1/genblk1[3].mult/added[1] ), .Y(n10902) );
  INVX1 U7639 ( .A(n11411), .Y(n10903) );
  NOR2X1 U7640 ( .A(n10903), .B(n10904), .Y(n10901) );
  NOR2X1 U7641 ( .A(n11412), .B(n10902), .Y(n10905) );
  INVX1 U7642 ( .A(n10905), .Y(n10904) );
  AND2X1 U7643 ( .A(n12147), .B(n12146), .Y(n12148) );
  INVX1 U7644 ( .A(n12148), .Y(n10906) );
  AND2X1 U7645 ( .A(n12042), .B(n12041), .Y(n12043) );
  INVX1 U7646 ( .A(n12043), .Y(n10907) );
  AND2X1 U7647 ( .A(n12077), .B(n12076), .Y(n12078) );
  INVX1 U7648 ( .A(n12078), .Y(n10908) );
  BUFX2 U7649 ( .A(n11501), .Y(n10909) );
  BUFX2 U7650 ( .A(n12794), .Y(n10910) );
  AND2X1 U7651 ( .A(\lamb/scale_ds1/genblk1[2].mult/added[1] ), .B(n11672), 
        .Y(n11673) );
  INVX1 U7652 ( .A(n11673), .Y(n10911) );
  BUFX2 U7653 ( .A(n12737), .Y(n10912) );
  NAND2X1 U7654 ( .A(n10913), .B(n10914), .Y(n12737) );
  INVX1 U7655 ( .A(n12749), .Y(n10915) );
  INVX1 U7656 ( .A(n12739), .Y(n10916) );
  NAND2X1 U7657 ( .A(n12732), .B(n10915), .Y(n10913) );
  NAND2X1 U7658 ( .A(n12732), .B(n10916), .Y(n10914) );
  BUFX2 U7659 ( .A(n12352), .Y(n10917) );
  INVX1 U7660 ( .A(n10918), .Y(n13571) );
  INVX1 U7661 ( .A(n13568), .Y(n10919) );
  INVX1 U7662 ( .A(n10647), .Y(n10920) );
  NOR2X1 U7663 ( .A(n10920), .B(n10921), .Y(n10918) );
  NOR2X1 U7664 ( .A(n10919), .B(n13640), .Y(n10922) );
  INVX1 U7665 ( .A(n10922), .Y(n10921) );
  BUFX2 U7666 ( .A(n12403), .Y(n10923) );
  AND2X1 U7667 ( .A(n12400), .B(n12171), .Y(n12417) );
  AND2X1 U7668 ( .A(n12227), .B(n12228), .Y(n12229) );
  INVX1 U7669 ( .A(n12229), .Y(n10924) );
  BUFX2 U7670 ( .A(n12540), .Y(n10925) );
  OR2X1 U7671 ( .A(n11751), .B(n11743), .Y(n11744) );
  INVX1 U7672 ( .A(n11744), .Y(n10926) );
  AND2X1 U7673 ( .A(n11473), .B(n11523), .Y(n11483) );
  INVX1 U7674 ( .A(n11483), .Y(n10927) );
  INVX1 U7675 ( .A(n10928), .Y(n12494) );
  INVX1 U7676 ( .A(n12492), .Y(n10929) );
  INVX1 U7677 ( .A(n12493), .Y(n10930) );
  NOR2X1 U7678 ( .A(n10930), .B(n10931), .Y(n10928) );
  NOR2X1 U7679 ( .A(n10929), .B(n12491), .Y(n10932) );
  INVX1 U7680 ( .A(n10932), .Y(n10931) );
  BUFX2 U7681 ( .A(n11872), .Y(n10933) );
  INVX1 U7682 ( .A(n10934), .Y(n11522) );
  INVX1 U7683 ( .A(n11515), .Y(n10935) );
  INVX1 U7684 ( .A(n11516), .Y(n10936) );
  NOR2X1 U7685 ( .A(n10814), .B(n10937), .Y(n10934) );
  NOR2X1 U7686 ( .A(n10935), .B(n10936), .Y(n10938) );
  INVX1 U7687 ( .A(n10938), .Y(n10937) );
  BUFX2 U7688 ( .A(n11380), .Y(n10939) );
  AND2X1 U7689 ( .A(\lamb/scale_ds1/genblk1[3].mult/added[4] ), .B(n11301), 
        .Y(n11303) );
  INVX1 U7690 ( .A(n11303), .Y(n10940) );
  OR2X1 U7691 ( .A(n13206), .B(n13205), .Y(n13207) );
  INVX1 U7692 ( .A(n13207), .Y(n10941) );
  OR2X1 U7693 ( .A(n11923), .B(\lamb/scale_bs3/genblk1[0].mult/added[1] ), .Y(
        n11924) );
  INVX1 U7694 ( .A(n11924), .Y(n10942) );
  AND2X1 U7695 ( .A(n13867), .B(n13123), .Y(n13124) );
  INVX1 U7696 ( .A(n13124), .Y(n10943) );
  INVX1 U7697 ( .A(n10944), .Y(n11738) );
  INVX1 U7698 ( .A(n11737), .Y(n10945) );
  INVX1 U7699 ( .A(n11765), .Y(n10946) );
  INVX1 U7700 ( .A(n11757), .Y(n10947) );
  NOR2X1 U7701 ( .A(n10947), .B(n10948), .Y(n10944) );
  NOR2X1 U7702 ( .A(n10945), .B(n10946), .Y(n10949) );
  INVX1 U7703 ( .A(n10949), .Y(n10948) );
  AND2X1 U7704 ( .A(n12362), .B(n12361), .Y(n12363) );
  INVX1 U7705 ( .A(n12363), .Y(n10950) );
  INVX1 U7706 ( .A(n10951), .Y(n11566) );
  INVX1 U7707 ( .A(n11564), .Y(n10952) );
  INVX1 U7708 ( .A(n11565), .Y(n10953) );
  INVX1 U7709 ( .A(n11583), .Y(n10954) );
  NOR2X1 U7710 ( .A(n10954), .B(n10955), .Y(n10951) );
  NOR2X1 U7711 ( .A(n10952), .B(n10953), .Y(n10956) );
  INVX1 U7712 ( .A(n10956), .Y(n10955) );
  AND2X1 U7713 ( .A(n12664), .B(n12671), .Y(n12660) );
  INVX1 U7714 ( .A(n12660), .Y(n10957) );
  AND2X1 U7715 ( .A(n13643), .B(n13660), .Y(n13661) );
  AND2X1 U7716 ( .A(n11427), .B(n11426), .Y(n11428) );
  INVX1 U7717 ( .A(n11428), .Y(n10958) );
  INVX1 U7718 ( .A(n10959), .Y(n12244) );
  INVX1 U7719 ( .A(n12255), .Y(n10960) );
  INVX1 U7720 ( .A(n12267), .Y(n10961) );
  NOR2X1 U7721 ( .A(n10961), .B(n10962), .Y(n10959) );
  NOR2X1 U7722 ( .A(n10960), .B(n12181), .Y(n10963) );
  INVX1 U7723 ( .A(n10963), .Y(n10962) );
  AND2X1 U7724 ( .A(n10519), .B(n12242), .Y(n12267) );
  AND2X1 U7725 ( .A(n11359), .B(n11330), .Y(n11324) );
  INVX1 U7726 ( .A(n11324), .Y(n10964) );
  AND2X1 U7727 ( .A(n11621), .B(n11560), .Y(n11561) );
  INVX1 U7728 ( .A(n11561), .Y(n10965) );
  OR2X1 U7729 ( .A(n13064), .B(n13062), .Y(n13056) );
  INVX1 U7730 ( .A(n13056), .Y(n10966) );
  BUFX2 U7731 ( .A(n13838), .Y(n10967) );
  INVX1 U7732 ( .A(n12868), .Y(n10968) );
  BUFX2 U7733 ( .A(n11783), .Y(n10969) );
  AND2X1 U7734 ( .A(n11768), .B(n11767), .Y(n11769) );
  INVX1 U7735 ( .A(n11769), .Y(n10970) );
  AND2X1 U7736 ( .A(n10528), .B(n11394), .Y(n11395) );
  INVX1 U7737 ( .A(n11395), .Y(n10971) );
  AND2X1 U7738 ( .A(n11704), .B(n11703), .Y(n11705) );
  INVX1 U7739 ( .A(n11705), .Y(n10972) );
  AND2X1 U7740 ( .A(n12335), .B(n12334), .Y(n12336) );
  INVX1 U7741 ( .A(n12336), .Y(n10973) );
  BUFX2 U7742 ( .A(n13774), .Y(n10974) );
  NOR2X1 U7743 ( .A(n10975), .B(n10976), .Y(n13774) );
  INVX1 U7744 ( .A(n13818), .Y(n10977) );
  NOR2X1 U7745 ( .A(n10977), .B(n13773), .Y(n10975) );
  INVX1 U7746 ( .A(n13816), .Y(n10978) );
  NOR2X1 U7747 ( .A(n10978), .B(n13772), .Y(n10976) );
  AND2X1 U7748 ( .A(n11862), .B(n11878), .Y(n11875) );
  INVX1 U7749 ( .A(n11875), .Y(n10979) );
  AND2X1 U7750 ( .A(n10675), .B(n11988), .Y(n11998) );
  INVX1 U7751 ( .A(n11998), .Y(n10980) );
  BUFX2 U7752 ( .A(\forney/m0/logB [3]), .Y(n10981) );
  AND2X1 U7753 ( .A(n11165), .B(n12957), .Y(n12959) );
  BUFX2 U7754 ( .A(n12619), .Y(n10982) );
  AND2X1 U7755 ( .A(n12564), .B(n12563), .Y(n12565) );
  INVX1 U7756 ( .A(n12565), .Y(n10983) );
  AND2X1 U7757 ( .A(n13893), .B(n12797), .Y(n12799) );
  INVX1 U7758 ( .A(n12799), .Y(n10984) );
  AND2X1 U7759 ( .A(n12558), .B(n12557), .Y(n12603) );
  INVX1 U7760 ( .A(n12603), .Y(n10985) );
  AND2X1 U7761 ( .A(n13590), .B(n12852), .Y(n12961) );
  INVX1 U7762 ( .A(n12961), .Y(n10986) );
  AND2X1 U7763 ( .A(\lamb/scale_ds1/genblk1[1].mult/added[3] ), .B(n12328), 
        .Y(n12310) );
  INVX1 U7764 ( .A(n12310), .Y(n10987) );
  AND2X1 U7765 ( .A(\add_x_135/n1 ), .B(
        \lamb/scale_ds2/genblk1[1].mult/added[4] ), .Y(n12217) );
  INVX1 U7766 ( .A(n12217), .Y(n10988) );
  INVX1 U7767 ( .A(n12988), .Y(n10989) );
  AND2X1 U7768 ( .A(n10621), .B(n11491), .Y(n11504) );
  INVX1 U7769 ( .A(n11504), .Y(n10990) );
  BUFX2 U7770 ( .A(n13407), .Y(n10991) );
  AND2X1 U7771 ( .A(n10644), .B(n13396), .Y(n13413) );
  AND2X1 U7772 ( .A(n13901), .B(n10477), .Y(n12934) );
  INVX1 U7773 ( .A(n12934), .Y(n10992) );
  AND2X1 U7774 ( .A(n12462), .B(n12440), .Y(n12461) );
  INVX1 U7775 ( .A(n12461), .Y(n10993) );
  OR2X1 U7776 ( .A(n12439), .B(n12460), .Y(n12462) );
  BUFX2 U7777 ( .A(n11451), .Y(n10994) );
  AND2X1 U7778 ( .A(n13160), .B(n13157), .Y(n13159) );
  INVX1 U7779 ( .A(n13159), .Y(n10995) );
  AND2X1 U7780 ( .A(n13069), .B(n13070), .Y(n13079) );
  INVX1 U7781 ( .A(n13079), .Y(n10996) );
  AND2X1 U7782 ( .A(n13065), .B(n10996), .Y(n13066) );
  BUFX2 U7783 ( .A(n11559), .Y(n10997) );
  AND2X1 U7784 ( .A(n10456), .B(n13457), .Y(n13471) );
  INVX1 U7785 ( .A(n13471), .Y(n10998) );
  AND2X1 U7786 ( .A(n12319), .B(\lamb/scale_ts1/genblk1[1].mult/added[1] ), 
        .Y(n12343) );
  INVX1 U7787 ( .A(n12343), .Y(n10999) );
  AND2X1 U7788 ( .A(n12240), .B(n12256), .Y(n12264) );
  INVX1 U7789 ( .A(n12264), .Y(n11000) );
  AND2X1 U7790 ( .A(\lamb/scale_ls2/genblk1[1].mult/added[2] ), .B(
        \lamb/scale_ls2/genblk1[1].mult/added[1] ), .Y(n11834) );
  INVX1 U7791 ( .A(n11834), .Y(n11001) );
  AND2X1 U7792 ( .A(\lamb/scale_ts2/genblk1[3].mult/added[1] ), .B(n11725), 
        .Y(n11730) );
  INVX1 U7793 ( .A(n11730), .Y(n11002) );
  BUFX2 U7794 ( .A(n12751), .Y(n11003) );
  BUFX2 U7795 ( .A(n11901), .Y(n11004) );
  NAND2X1 U7796 ( .A(n11005), .B(n11006), .Y(n11901) );
  INVX1 U7797 ( .A(n11816), .Y(n11007) );
  INVX1 U7798 ( .A(n10507), .Y(n11008) );
  NAND2X1 U7799 ( .A(n11957), .B(n11007), .Y(n11005) );
  NAND2X1 U7800 ( .A(n11957), .B(n11008), .Y(n11006) );
  INVX1 U7801 ( .A(n11009), .Y(n13259) );
  INVX1 U7802 ( .A(n11709), .Y(n11010) );
  NOR2X1 U7803 ( .A(n11711), .B(n11011), .Y(n11009) );
  NOR2X1 U7804 ( .A(n12678), .B(n11010), .Y(n11012) );
  INVX1 U7805 ( .A(n11012), .Y(n11011) );
  INVX1 U7806 ( .A(n12498), .Y(n11013) );
  BUFX2 U7807 ( .A(n13404), .Y(n11014) );
  AND2X1 U7808 ( .A(n10849), .B(n12706), .Y(n12701) );
  INVX1 U7809 ( .A(n12701), .Y(n11015) );
  AND2X1 U7810 ( .A(n12219), .B(n12221), .Y(n12253) );
  INVX1 U7811 ( .A(n12253), .Y(n11016) );
  AND2X1 U7812 ( .A(n13545), .B(n13544), .Y(n13558) );
  INVX1 U7813 ( .A(n13558), .Y(n11017) );
  BUFX2 U7814 ( .A(n12381), .Y(n11018) );
  AND2X1 U7815 ( .A(n13011), .B(n12633), .Y(n12628) );
  INVX1 U7816 ( .A(n12628), .Y(n11019) );
  INVX1 U7817 ( .A(n13264), .Y(n11020) );
  AND2X1 U7818 ( .A(\lamb/scale_ds2/genblk1[1].mult/added[2] ), .B(n12230), 
        .Y(n12249) );
  INVX1 U7819 ( .A(n12249), .Y(n11021) );
  AND2X1 U7820 ( .A(n12294), .B(n10618), .Y(n12302) );
  INVX1 U7821 ( .A(n12302), .Y(n11022) );
  BUFX2 U7822 ( .A(n13155), .Y(n11023) );
  AND2X1 U7823 ( .A(n11314), .B(n12680), .Y(n13382) );
  INVX1 U7824 ( .A(n13382), .Y(n11024) );
  BUFX2 U7825 ( .A(n12942), .Y(n11025) );
  INVX1 U7826 ( .A(n11026), .Y(n12394) );
  INVX1 U7827 ( .A(n12284), .Y(n11027) );
  INVX1 U7828 ( .A(n12285), .Y(n11028) );
  NOR2X1 U7829 ( .A(n10682), .B(n11029), .Y(n11026) );
  NOR2X1 U7830 ( .A(n11027), .B(n11028), .Y(n11030) );
  INVX1 U7831 ( .A(n11030), .Y(n11029) );
  AND2X1 U7832 ( .A(n12511), .B(n13154), .Y(n13163) );
  INVX1 U7833 ( .A(n13163), .Y(n11031) );
  AND2X1 U7834 ( .A(n11031), .B(n13168), .Y(n13151) );
  INVX1 U7835 ( .A(n10364), .Y(n11032) );
  BUFX2 U7836 ( .A(\lamb/scale_ts3/genblk1[3].mult/logA[2] ), .Y(n11033) );
  NAND2X1 U7837 ( .A(n11034), .B(n11035), .Y(
        \lamb/scale_ts3/genblk1[3].mult/logA[2] ) );
  INVX1 U7838 ( .A(n13029), .Y(n11036) );
  INVX1 U7839 ( .A(n13033), .Y(n11037) );
  INVX1 U7840 ( .A(n10543), .Y(n11038) );
  NAND2X1 U7841 ( .A(n11036), .B(n11037), .Y(n11034) );
  NAND2X1 U7842 ( .A(n11036), .B(n11038), .Y(n11035) );
  BUFX2 U7843 ( .A(\lamb/scale_ts3/genblk1[2].mult/logA[2] ), .Y(n11039) );
  INVX1 U7844 ( .A(n11040), .Y(n10368) );
  INVX1 U7845 ( .A(n13870), .Y(n11041) );
  INVX1 U7846 ( .A(n13871), .Y(n11042) );
  INVX1 U7847 ( .A(n10549), .Y(n11043) );
  NOR2X1 U7848 ( .A(n11043), .B(n11044), .Y(n11040) );
  NOR2X1 U7849 ( .A(n11041), .B(n11042), .Y(n11045) );
  INVX1 U7850 ( .A(n11045), .Y(n11044) );
  OR2X1 U7851 ( .A(n10817), .B(n10492), .Y(n13871) );
  BUFX2 U7852 ( .A(\lamb/scale_ts2/genblk1[2].mult/logA[2] ), .Y(n11046) );
  BUFX2 U7853 ( .A(\lamb/scale_ts0/genblk1[1].mult/logA[2] ), .Y(n11047) );
  AND2X1 U7854 ( .A(n11503), .B(n11484), .Y(n11489) );
  INVX1 U7855 ( .A(n11489), .Y(n11048) );
  INVX1 U7856 ( .A(n12847), .Y(n11049) );
  AND2X1 U7857 ( .A(n10552), .B(n11419), .Y(n11444) );
  INVX1 U7858 ( .A(n11444), .Y(n11050) );
  BUFX2 U7859 ( .A(n11802), .Y(n11051) );
  AND2X1 U7860 ( .A(n11299), .B(n11298), .Y(n11440) );
  INVX1 U7861 ( .A(n11440), .Y(n11052) );
  BUFX2 U7862 ( .A(n12340), .Y(n11053) );
  AND2X1 U7863 ( .A(n13194), .B(n13879), .Y(n13882) );
  INVX1 U7864 ( .A(n13882), .Y(n11054) );
  BUFX2 U7865 ( .A(n12872), .Y(n11055) );
  AND2X1 U7866 ( .A(n10831), .B(n13943), .Y(n13185) );
  INVX1 U7867 ( .A(n13185), .Y(n11056) );
  AND2X1 U7868 ( .A(n12298), .B(n12297), .Y(n12358) );
  INVX1 U7869 ( .A(n12358), .Y(n11057) );
  AND2X1 U7870 ( .A(n13274), .B(n13269), .Y(n13278) );
  INVX1 U7871 ( .A(n13278), .Y(n11058) );
  AND2X1 U7872 ( .A(n12428), .B(n12536), .Y(n12576) );
  INVX1 U7873 ( .A(n12576), .Y(n11059) );
  BUFX2 U7874 ( .A(n12925), .Y(n11060) );
  INVX1 U7875 ( .A(n11061), .Y(n12755) );
  INVX1 U7876 ( .A(n10513), .Y(n11062) );
  INVX1 U7877 ( .A(n12741), .Y(n11063) );
  NOR2X1 U7878 ( .A(n11063), .B(n11064), .Y(n11061) );
  NOR2X1 U7879 ( .A(\lamb/scale_ts1/genblk1[0].mult/added[1] ), .B(n11062), 
        .Y(n11065) );
  INVX1 U7880 ( .A(n11065), .Y(n11064) );
  INVX1 U7881 ( .A(n11066), .Y(n11885) );
  INVX1 U7882 ( .A(n11863), .Y(n11067) );
  INVX1 U7883 ( .A(n11864), .Y(n11068) );
  NOR2X1 U7884 ( .A(n11068), .B(n11069), .Y(n11066) );
  NOR2X1 U7885 ( .A(n10731), .B(n11067), .Y(n11070) );
  INVX1 U7886 ( .A(n11070), .Y(n11069) );
  BUFX2 U7887 ( .A(n13293), .Y(n11071) );
  NOR2X1 U7888 ( .A(n11072), .B(n11073), .Y(n13293) );
  INVX1 U7889 ( .A(n11075), .Y(n11074) );
  NOR2X1 U7890 ( .A(n10795), .B(n11074), .Y(n11072) );
  INVX1 U7891 ( .A(n13280), .Y(n11075) );
  NOR2X1 U7892 ( .A(n11075), .B(n10794), .Y(n11073) );
  OR2X1 U7893 ( .A(n13099), .B(n13100), .Y(n13096) );
  INVX1 U7894 ( .A(n13096), .Y(n11076) );
  BUFX2 U7895 ( .A(n11601), .Y(n11077) );
  AND2X1 U7896 ( .A(n13342), .B(n13348), .Y(n13351) );
  INVX1 U7897 ( .A(n13351), .Y(n11078) );
  AND2X1 U7898 ( .A(n12807), .B(n12832), .Y(n12168) );
  INVX1 U7899 ( .A(n12168), .Y(n11079) );
  AND2X1 U7900 ( .A(n11661), .B(n11660), .Y(n11670) );
  INVX1 U7901 ( .A(n11670), .Y(n11080) );
  BUFX2 U7902 ( .A(n12582), .Y(n11081) );
  AND2X1 U7903 ( .A(n11546), .B(n11548), .Y(n11551) );
  INVX1 U7904 ( .A(n11551), .Y(n11082) );
  BUFX2 U7905 ( .A(n11690), .Y(n11083) );
  OR2X1 U7906 ( .A(n12989), .B(n12981), .Y(n12987) );
  INVX1 U7907 ( .A(n12987), .Y(n11084) );
  BUFX2 U7908 ( .A(n11507), .Y(n11085) );
  INVX1 U7909 ( .A(n11855), .Y(n11086) );
  AND2X1 U7910 ( .A(n12391), .B(n12390), .Y(n12410) );
  INVX1 U7911 ( .A(n12410), .Y(n11087) );
  INVX1 U7912 ( .A(n11088), .Y(n12502) );
  INVX1 U7913 ( .A(n12470), .Y(n11089) );
  INVX1 U7914 ( .A(n12471), .Y(n11090) );
  INVX1 U7915 ( .A(\lamb/scale_ds2/genblk1[2].mult/added[1] ), .Y(n11091) );
  NOR2X1 U7916 ( .A(n11091), .B(n11092), .Y(n11088) );
  NOR2X1 U7917 ( .A(n11089), .B(n11090), .Y(n11093) );
  INVX1 U7918 ( .A(n11093), .Y(n11092) );
  BUFX2 U7919 ( .A(n11268), .Y(n11094) );
  AND2X1 U7920 ( .A(n13053), .B(n13052), .Y(n13059) );
  INVX1 U7921 ( .A(n13059), .Y(n11095) );
  BUFX2 U7922 ( .A(n11259), .Y(n11096) );
  AND2X1 U7923 ( .A(n13640), .B(n13615), .Y(n13638) );
  INVX1 U7924 ( .A(n13638), .Y(n11097) );
  AND2X1 U7925 ( .A(\add_x_121/n1 ), .B(
        \lamb/scale_ds3/genblk1[2].mult/added[4] ), .Y(n12178) );
  INVX1 U7926 ( .A(n12178), .Y(n11098) );
  BUFX2 U7927 ( .A(n12396), .Y(n11099) );
  INVX1 U7928 ( .A(n11100), .Y(n11750) );
  INVX1 U7929 ( .A(n10510), .Y(n11101) );
  INVX1 U7930 ( .A(n11717), .Y(n11102) );
  NOR2X1 U7931 ( .A(n11102), .B(n11103), .Y(n11100) );
  NOR2X1 U7932 ( .A(n11101), .B(\lamb/scale_ts2/genblk1[3].mult/added[3] ), 
        .Y(n11104) );
  INVX1 U7933 ( .A(n11104), .Y(n11103) );
  BUFX2 U7934 ( .A(n11592), .Y(n11105) );
  OR2X1 U7935 ( .A(n11296), .B(n11302), .Y(n11300) );
  INVX1 U7936 ( .A(n11300), .Y(n11106) );
  BUFX2 U7937 ( .A(n11518), .Y(n11107) );
  AND2X1 U7938 ( .A(n10624), .B(n13527), .Y(n13551) );
  INVX1 U7939 ( .A(n13551), .Y(n11108) );
  INVX1 U7940 ( .A(n11109), .Y(n13924) );
  INVX1 U7941 ( .A(n12196), .Y(n11110) );
  INVX1 U7942 ( .A(n12195), .Y(n11111) );
  NOR2X1 U7943 ( .A(n12193), .B(n11112), .Y(n11109) );
  NOR2X1 U7944 ( .A(n11110), .B(n11111), .Y(n11113) );
  INVX1 U7945 ( .A(n11113), .Y(n11112) );
  AND2X1 U7946 ( .A(\lamb/scale_bs3/genblk1[0].mult/added[3] ), .B(n11806), 
        .Y(n11927) );
  INVX1 U7947 ( .A(n11927), .Y(n11114) );
  INVX1 U7948 ( .A(n11453), .Y(n11115) );
  INVX1 U7949 ( .A(n12270), .Y(n11116) );
  AND2X1 U7950 ( .A(n13831), .B(n13332), .Y(n13828) );
  INVX1 U7951 ( .A(n13828), .Y(n11117) );
  AND2X1 U7952 ( .A(n11117), .B(n10498), .Y(n13829) );
  AND2X1 U7953 ( .A(n13350), .B(n13349), .Y(n13345) );
  INVX1 U7954 ( .A(n13345), .Y(n11118) );
  XOR2X1 U7955 ( .A(n11599), .B(n12667), .Y(n13349) );
  BUFX2 U7956 ( .A(n13356), .Y(n11119) );
  AND2X1 U7957 ( .A(n12916), .B(n10854), .Y(n12910) );
  INVX1 U7958 ( .A(n12910), .Y(n11120) );
  AND2X1 U7959 ( .A(n13193), .B(n13876), .Y(n13878) );
  INVX1 U7960 ( .A(n13878), .Y(n11121) );
  INVX1 U7961 ( .A(n11789), .Y(n11122) );
  INVX1 U7962 ( .A(n11310), .Y(n11123) );
  AND2X1 U7963 ( .A(n11293), .B(n11292), .Y(n13255) );
  INVX1 U7964 ( .A(n13255), .Y(n11124) );
  AND2X1 U7965 ( .A(n13140), .B(n13141), .Y(n13148) );
  INVX1 U7966 ( .A(n13148), .Y(n11125) );
  AND2X1 U7967 ( .A(\lamb/scale_ls2/genblk1[2].mult/added[4] ), .B(
        \add_x_139/n1 ), .Y(n13106) );
  INVX1 U7968 ( .A(n13106), .Y(n11126) );
  AND2X1 U7969 ( .A(n12293), .B(n13370), .Y(n13824) );
  INVX1 U7970 ( .A(n13824), .Y(n11127) );
  AND2X1 U7971 ( .A(n11637), .B(n11636), .Y(n11695) );
  INVX1 U7972 ( .A(n11695), .Y(n11128) );
  INVX1 U7973 ( .A(n12922), .Y(n11129) );
  INVX1 U7974 ( .A(n12545), .Y(n11130) );
  AND2X1 U7975 ( .A(\add_x_128/n1 ), .B(
        \lamb/scale_ls3/genblk1[0].mult/added[4] ), .Y(n11542) );
  INVX1 U7976 ( .A(n11542), .Y(n11131) );
  AND2X1 U7977 ( .A(\forney/pe0/mult0/added [4]), .B(\add_x_87/n1 ), .Y(n12572) );
  INVX1 U7978 ( .A(n12572), .Y(n11132) );
  AND2X1 U7979 ( .A(n12665), .B(n12667), .Y(n12668) );
  INVX1 U7980 ( .A(n12668), .Y(n11133) );
  AND2X1 U7981 ( .A(n13354), .B(n13927), .Y(n13362) );
  INVX1 U7982 ( .A(n13362), .Y(n11134) );
  INVX1 U7983 ( .A(n12970), .Y(n11135) );
  OR2X1 U7984 ( .A(n13108), .B(n10673), .Y(n13113) );
  INVX1 U7985 ( .A(n13113), .Y(n11136) );
  AND2X1 U7986 ( .A(n13834), .B(n13337), .Y(n13833) );
  INVX1 U7987 ( .A(n13833), .Y(n11137) );
  OR2X1 U7988 ( .A(n13122), .B(n13121), .Y(n13866) );
  INVX1 U7989 ( .A(n13866), .Y(n11138) );
  OR2X1 U7990 ( .A(n13935), .B(n13933), .Y(n13941) );
  INVX1 U7991 ( .A(n13941), .Y(n11139) );
  AND2X1 U7992 ( .A(n10540), .B(n13531), .Y(n13539) );
  INVX1 U7993 ( .A(n13539), .Y(n11140) );
  AND2X1 U7994 ( .A(\forney/m0/added [3]), .B(n13389), .Y(n13391) );
  INVX1 U7995 ( .A(n13391), .Y(n11141) );
  BUFX2 U7996 ( .A(n13649), .Y(n11142) );
  AND2X1 U7997 ( .A(\lamb/scale_ls3/genblk1[1].mult/added[1] ), .B(
        \lamb/scale_ls3/genblk1[1].mult/added[2] ), .Y(n11963) );
  INVX1 U7998 ( .A(n11963), .Y(n11143) );
  OR2X1 U7999 ( .A(\lamb/scale_ds1/genblk1[3].mult/added[3] ), .B(n11430), .Y(
        n11457) );
  INVX1 U8000 ( .A(n11457), .Y(n11144) );
  BUFX2 U8001 ( .A(n12642), .Y(n11145) );
  AND2X1 U8002 ( .A(n13058), .B(n13057), .Y(n12616) );
  INVX1 U8003 ( .A(n12616), .Y(n11146) );
  BUFX2 U8004 ( .A(n12356), .Y(n11147) );
  BUFX2 U8005 ( .A(n12602), .Y(n11148) );
  AND2X1 U8006 ( .A(n13001), .B(n12630), .Y(n13002) );
  BUFX2 U8007 ( .A(n12495), .Y(n11149) );
  BUFX2 U8008 ( .A(n13308), .Y(n11150) );
  AND2X1 U8009 ( .A(\lamb/scale_ds2/genblk1[3].mult/added[4] ), .B(
        \add_x_133/n1 ), .Y(n11759) );
  INVX1 U8010 ( .A(n11759), .Y(n11151) );
  BUFX2 U8011 ( .A(n11459), .Y(n11152) );
  AND2X1 U8012 ( .A(n13341), .B(n13340), .Y(n11693) );
  INVX1 U8013 ( .A(n11693), .Y(n11153) );
  AND2X1 U8014 ( .A(n13201), .B(n13202), .Y(n12505) );
  INVX1 U8015 ( .A(n12505), .Y(n11154) );
  AND2X1 U8016 ( .A(n13067), .B(n13076), .Y(n12422) );
  INVX1 U8017 ( .A(n12422), .Y(n11155) );
  BUFX2 U8018 ( .A(n11626), .Y(n11156) );
  AND2X1 U8019 ( .A(n13693), .B(n13387), .Y(n12620) );
  INVX1 U8020 ( .A(n12620), .Y(n11157) );
  OR2X1 U8021 ( .A(n10585), .B(n13458), .Y(n13547) );
  INVX1 U8022 ( .A(n13547), .Y(n11158) );
  BUFX2 U8023 ( .A(n11505), .Y(n11159) );
  BUFX2 U8024 ( .A(n11349), .Y(n11160) );
  BUFX2 U8025 ( .A(n12849), .Y(n11161) );
  OR2X1 U8026 ( .A(n10447), .B(n11161), .Y(n12855) );
  BUFX2 U8027 ( .A(n13538), .Y(n11162) );
  OR2X1 U8028 ( .A(n13455), .B(n11162), .Y(n13463) );
  OR2X1 U8029 ( .A(n12974), .B(n13487), .Y(n12997) );
  INVX1 U8030 ( .A(n12997), .Y(n11163) );
  AND2X1 U8031 ( .A(n13602), .B(n10612), .Y(n13003) );
  INVX1 U8032 ( .A(n13003), .Y(n11164) );
  AND2X1 U8033 ( .A(n12952), .B(n12951), .Y(n12956) );
  INVX1 U8034 ( .A(n12956), .Y(n11165) );
  AND2X1 U8035 ( .A(n11650), .B(n11676), .Y(n11688) );
  INVX1 U8036 ( .A(n11688), .Y(n11166) );
  BUFX2 U8037 ( .A(n12652), .Y(n11167) );
  INVX1 U8038 ( .A(n11761), .Y(n11168) );
  BUFX2 U8039 ( .A(n13242), .Y(n11169) );
  AND2X1 U8040 ( .A(n13662), .B(n13623), .Y(n13706) );
  INVX1 U8041 ( .A(n13706), .Y(n11170) );
  AND2X1 U8042 ( .A(n13667), .B(n13684), .Y(n13674) );
  INVX1 U8043 ( .A(n13674), .Y(n11171) );
  AND2X1 U8044 ( .A(n13489), .B(n12804), .Y(n13582) );
  INVX1 U8045 ( .A(n13582), .Y(n11172) );
  OR2X1 U8046 ( .A(\lamb/scale_ts0/genblk1[2].mult/added[4] ), .B(
        \add_x_152/n1 ), .Y(n11329) );
  INVX1 U8047 ( .A(n11329), .Y(n11173) );
  AND2X1 U8048 ( .A(n13229), .B(n12760), .Y(n13230) );
  INVX1 U8049 ( .A(n13230), .Y(n11174) );
  BUFX2 U8050 ( .A(n13749), .Y(n11175) );
  AND2X1 U8051 ( .A(n13602), .B(n13598), .Y(n13599) );
  AND2X1 U8052 ( .A(n10567), .B(n12983), .Y(n12990) );
  INVX1 U8053 ( .A(n12990), .Y(n11176) );
  AND2X1 U8054 ( .A(n12767), .B(n13143), .Y(n13142) );
  INVX1 U8055 ( .A(n13142), .Y(n11177) );
  BUFX2 U8056 ( .A(\forney/pe0/mult0/logA [2]), .Y(n11178) );
  INVX1 U8057 ( .A(n11179), .Y(n13542) );
  NAND2X1 U8058 ( .A(n13520), .B(n13519), .Y(n11180) );
  NAND2X1 U8059 ( .A(n13518), .B(n13517), .Y(n11181) );
  NAND2X1 U8060 ( .A(n11180), .B(n11181), .Y(n11179) );
  INVX1 U8061 ( .A(n12387), .Y(n11182) );
  AND2X1 U8062 ( .A(\add_x_148/n1 ), .B(
        \lamb/scale_ds1/genblk1[1].mult/added[4] ), .Y(n12330) );
  INVX1 U8063 ( .A(n12330), .Y(n11183) );
  AND2X1 U8064 ( .A(\lamb/scale_ts0/genblk1[0].mult/added[3] ), .B(n12186), 
        .Y(n12209) );
  INVX1 U8065 ( .A(n12209), .Y(n11184) );
  INVX1 U8066 ( .A(n11185), .Y(n13917) );
  INVX1 U8067 ( .A(n12746), .Y(n11186) );
  INVX1 U8068 ( .A(n12747), .Y(n11187) );
  INVX1 U8069 ( .A(n12752), .Y(n11188) );
  NOR2X1 U8070 ( .A(n11188), .B(n11189), .Y(n11185) );
  NOR2X1 U8071 ( .A(n11186), .B(n11187), .Y(n11190) );
  INVX1 U8072 ( .A(n11190), .Y(n11189) );
  BUFX2 U8073 ( .A(n11368), .Y(n11191) );
  AND2X1 U8074 ( .A(n13586), .B(n12935), .Y(n12858) );
  INVX1 U8075 ( .A(n12858), .Y(n11192) );
  AND2X1 U8076 ( .A(\lamb/scale_ds3/genblk1[3].mult/added[2] ), .B(
        \lamb/scale_ds3/genblk1[3].mult/added[1] ), .Y(n12549) );
  INVX1 U8077 ( .A(n12549), .Y(n11193) );
  AND2X1 U8078 ( .A(\lamb/scale_ls3/genblk1[2].mult/added[4] ), .B(
        \add_x_126/n1 ), .Y(n11937) );
  INVX1 U8079 ( .A(n11937), .Y(n11194) );
  AND2X1 U8080 ( .A(n10450), .B(n12833), .Y(n13691) );
  INVX1 U8081 ( .A(n13691), .Y(n11195) );
  AND2X1 U8082 ( .A(n13431), .B(n11909), .Y(n13442) );
  INVX1 U8083 ( .A(n13442), .Y(n11196) );
  OR2X1 U8084 ( .A(\forney/m1/added [4]), .B(\add_x_20/n1 ), .Y(n13513) );
  INVX1 U8085 ( .A(n13513), .Y(n11197) );
  AND2X1 U8086 ( .A(n12822), .B(n13903), .Y(n13695) );
  INVX1 U8087 ( .A(n13695), .Y(n11198) );
  INVX1 U8088 ( .A(n11199), .Y(n13267) );
  NAND2X1 U8089 ( .A(n10851), .B(n11712), .Y(n11200) );
  NAND2X1 U8090 ( .A(n13371), .B(n12682), .Y(n11201) );
  NAND2X1 U8091 ( .A(n11200), .B(n11201), .Y(n11199) );
  OR2X1 U8092 ( .A(n13411), .B(n13410), .Y(n13451) );
  INVX1 U8093 ( .A(n13451), .Y(n11202) );
  INVX1 U8094 ( .A(n13588), .Y(n11203) );
  BUFX2 U8095 ( .A(\lamb/scale_bs3/genblk1[0].mult/logB[3] ), .Y(n11204) );
  BUFX2 U8096 ( .A(\lamb/scale_bs2/genblk1[1].mult/added[4] ), .Y(n11205) );
  AND2X1 U8097 ( .A(n13847), .B(n13856), .Y(n13862) );
  BUFX2 U8098 ( .A(\lamb/scale_ts1/genblk1[0].mult/logB[3] ), .Y(n11206) );
  AND2X1 U8099 ( .A(\add_x_85/n1 ), .B(\forney/pe1/mult0/added [4]), .Y(n12881) );
  INVX1 U8100 ( .A(n12881), .Y(n11207) );
  BUFX2 U8101 ( .A(n13634), .Y(n11208) );
  INVX1 U8102 ( .A(n13218), .Y(n11209) );
  AND2X1 U8103 ( .A(n13896), .B(n12964), .Y(n13888) );
  INVX1 U8104 ( .A(n13888), .Y(n11210) );
  BUFX2 U8105 ( .A(\lamb/scale_bs3/genblk1[0].mult/logB[1] ), .Y(n11211) );
  BUFX2 U8106 ( .A(\lamb/scale_bs2/genblk1[1].mult/added[2] ), .Y(n11212) );
  BUFX2 U8107 ( .A(\lamb/scale_ts1/genblk1[0].mult/logB[1] ), .Y(n11213) );
  BUFX2 U8108 ( .A(\lamb/scale_ts1/genblk1[0].mult/logB[2] ), .Y(n11214) );
  NAND2X1 U8109 ( .A(n11215), .B(n11216), .Y(
        \lamb/scale_ts1/genblk1[0].mult/logB[2] ) );
  INVX1 U8110 ( .A(n13321), .Y(n11217) );
  INVX1 U8111 ( .A(n13322), .Y(n11218) );
  INVX1 U8112 ( .A(n13323), .Y(n11219) );
  NAND2X1 U8113 ( .A(n11217), .B(n11218), .Y(n11215) );
  NAND2X1 U8114 ( .A(n11217), .B(n11219), .Y(n11216) );
  INVX1 U8115 ( .A(n11220), .Y(n12132) );
  INVX1 U8116 ( .A(n11949), .Y(n11221) );
  INVX1 U8117 ( .A(n11950), .Y(n11222) );
  INVX1 U8118 ( .A(n11951), .Y(n11223) );
  NOR2X1 U8119 ( .A(n11223), .B(n11224), .Y(n11220) );
  NOR2X1 U8120 ( .A(n11221), .B(n11222), .Y(n11225) );
  INVX1 U8121 ( .A(n11225), .Y(n11224) );
  BUFX2 U8122 ( .A(\lamb/scale_ls3/genblk1[0].mult/logB[2] ), .Y(n11226) );
  BUFX2 U8123 ( .A(n13086), .Y(n11227) );
  OR2X1 U8124 ( .A(n13752), .B(n13751), .Y(n13686) );
  INVX1 U8125 ( .A(n13686), .Y(n11228) );
  OR2X1 U8126 ( .A(n13747), .B(n10753), .Y(n13741) );
  INVX1 U8127 ( .A(n13741), .Y(n11229) );
  BUFX2 U8128 ( .A(\lamb/scale_ls2/genblk1[0].mult/logB[2] ), .Y(n11230) );
  OR2X1 U8129 ( .A(n13228), .B(n12764), .Y(n10375) );
  INVX1 U8130 ( .A(n10375), .Y(n11231) );
  AND2X1 U8131 ( .A(n12695), .B(n11646), .Y(n13235) );
  INVX1 U8132 ( .A(msg[32]), .Y(n13688) );
  INVX1 U8133 ( .A(msg[24]), .Y(n13725) );
  INVX1 U8134 ( .A(msg[4]), .Y(n13803) );
  AOI22X1 U8135 ( .A(msg[4]), .B(msg[24]), .C(n13725), .D(n13803), .Y(n11592)
         );
  MUX2X1 U8136 ( .B(n13688), .A(msg[32]), .S(n11105), .Y(n11266) );
  INVX1 U8137 ( .A(msg[23]), .Y(n13727) );
  INVX1 U8138 ( .A(msg[26]), .Y(n13721) );
  AOI22X1 U8139 ( .A(msg[26]), .B(n13727), .C(msg[23]), .D(n13721), .Y(n11232)
         );
  INVX1 U8140 ( .A(n11232), .Y(n11591) );
  HAX1 U8141 ( .A(n11266), .B(n11591), .YS(n13311) );
  INVX1 U8142 ( .A(msg[52]), .Y(n11336) );
  INVX1 U8143 ( .A(msg[22]), .Y(n13729) );
  MUX2X1 U8144 ( .B(n13729), .A(msg[22]), .S(msg[46]), .Y(n11271) );
  MUX2X1 U8145 ( .B(n11336), .A(msg[52]), .S(n11271), .Y(n11364) );
  HAX1 U8146 ( .A(n13311), .B(n11364), .YS(n11577) );
  INVX1 U8147 ( .A(msg[18]), .Y(n13737) );
  INVX1 U8148 ( .A(msg[42]), .Y(n13625) );
  MUX2X1 U8149 ( .B(msg[42]), .A(n13625), .S(msg[58]), .Y(n12645) );
  INVX1 U8150 ( .A(msg[15]), .Y(n13758) );
  INVX1 U8151 ( .A(msg[48]), .Y(n12646) );
  AOI22X1 U8152 ( .A(msg[48]), .B(n13758), .C(msg[15]), .D(n12646), .Y(n11259)
         );
  HAX1 U8153 ( .A(n12645), .B(n11096), .YS(n11233) );
  MUX2X1 U8154 ( .B(n13737), .A(msg[18]), .S(n11233), .Y(n13312) );
  INVX1 U8155 ( .A(msg[28]), .Y(n13717) );
  INVX1 U8156 ( .A(msg[20]), .Y(n13733) );
  INVX1 U8157 ( .A(msg[40]), .Y(n13666) );
  MUX2X1 U8158 ( .B(msg[20]), .A(n13733), .S(n13666), .Y(n11254) );
  MUX2X1 U8159 ( .B(n13717), .A(msg[28]), .S(n11254), .Y(n11270) );
  INVX1 U8160 ( .A(msg[19]), .Y(n13735) );
  INVX1 U8161 ( .A(msg[39]), .Y(n13669) );
  MUX2X1 U8162 ( .B(msg[19]), .A(n13735), .S(n13669), .Y(n11288) );
  HAX1 U8163 ( .A(n11270), .B(n11288), .YS(n11234) );
  FAX1 U8164 ( .A(n11577), .B(n13312), .C(n11234), .YS(n11387) );
  INVX1 U8165 ( .A(msg[14]), .Y(n13761) );
  INVX1 U8166 ( .A(msg[34]), .Y(n13681) );
  MUX2X1 U8167 ( .B(msg[14]), .A(n13761), .S(n13681), .Y(n11384) );
  INVX1 U8168 ( .A(msg[31]), .Y(n13705) );
  INVX1 U8169 ( .A(msg[17]), .Y(n13739) );
  INVX1 U8170 ( .A(msg[37]), .Y(n13673) );
  MUX2X1 U8171 ( .B(msg[17]), .A(n13739), .S(n13673), .Y(n11369) );
  MUX2X1 U8172 ( .B(n13705), .A(msg[31]), .S(n11369), .Y(n11241) );
  HAX1 U8173 ( .A(n11384), .B(n11241), .YS(n11247) );
  INVX1 U8174 ( .A(msg[21]), .Y(n13731) );
  INVX1 U8175 ( .A(msg[29]), .Y(n13711) );
  INVX1 U8176 ( .A(msg[25]), .Y(n13723) );
  INVX1 U8177 ( .A(msg[45]), .Y(n11235) );
  AOI22X1 U8178 ( .A(msg[45]), .B(msg[25]), .C(n13723), .D(n11235), .Y(n12642)
         );
  INVX1 U8179 ( .A(n11145), .Y(n12641) );
  MUX2X1 U8180 ( .B(msg[29]), .A(n13711), .S(n12641), .Y(n11236) );
  MUX2X1 U8181 ( .B(n13731), .A(msg[21]), .S(n11236), .Y(n11238) );
  INVX1 U8182 ( .A(msg[1]), .Y(n13815) );
  INVX1 U8183 ( .A(msg[11]), .Y(n13775) );
  INVX1 U8184 ( .A(msg[43]), .Y(n13604) );
  MUX2X1 U8185 ( .B(n13604), .A(msg[43]), .S(msg[55]), .Y(n11392) );
  MUX2X1 U8186 ( .B(n13775), .A(msg[11]), .S(n11392), .Y(n11284) );
  MUX2X1 U8187 ( .B(n13815), .A(msg[1]), .S(n11284), .Y(n11237) );
  FAX1 U8188 ( .A(msg[49]), .B(n11238), .C(n11237), .YS(n11239) );
  FAX1 U8189 ( .A(n11387), .B(n11247), .C(n11239), .YS(n11712) );
  INVX1 U8190 ( .A(msg[59]), .Y(n13300) );
  INVX1 U8191 ( .A(msg[6]), .Y(n13795) );
  INVX1 U8192 ( .A(msg[3]), .Y(n13807) );
  MUX2X1 U8193 ( .B(msg[6]), .A(n13795), .S(n13807), .Y(n13298) );
  INVX1 U8194 ( .A(n13298), .Y(n13299) );
  MUX2X1 U8195 ( .B(n13604), .A(msg[43]), .S(n13299), .Y(n11570) );
  HAX1 U8196 ( .A(n11384), .B(n11570), .YS(n11337) );
  MUX2X1 U8197 ( .B(msg[59]), .A(n13300), .S(n11337), .Y(n11319) );
  INVX1 U8198 ( .A(msg[8]), .Y(n13787) );
  INVX1 U8199 ( .A(msg[36]), .Y(n13677) );
  AOI22X1 U8200 ( .A(msg[36]), .B(msg[8]), .C(n13787), .D(n13677), .Y(n11349)
         );
  INVX1 U8201 ( .A(msg[12]), .Y(n13770) );
  INVX1 U8202 ( .A(msg[16]), .Y(n13743) );
  MUX2X1 U8203 ( .B(msg[12]), .A(n13770), .S(n13743), .Y(n11249) );
  HAX1 U8204 ( .A(n11160), .B(n11249), .YS(n13306) );
  INVX1 U8205 ( .A(n13306), .Y(n13305) );
  INVX1 U8206 ( .A(msg[9]), .Y(n13783) );
  MUX2X1 U8207 ( .B(n13783), .A(msg[9]), .S(msg[49]), .Y(n11279) );
  HAX1 U8208 ( .A(n11254), .B(n11279), .YS(n11587) );
  INVX1 U8209 ( .A(n11587), .Y(n11240) );
  HAX1 U8210 ( .A(n13305), .B(n11240), .YS(n11339) );
  INVX1 U8211 ( .A(msg[7]), .Y(n13791) );
  INVX1 U8212 ( .A(msg[10]), .Y(n13779) );
  AOI22X1 U8213 ( .A(msg[10]), .B(msg[7]), .C(n13791), .D(n13779), .Y(n11368)
         );
  MUX2X1 U8214 ( .B(n13717), .A(msg[28]), .S(n11191), .Y(n11398) );
  INVX1 U8215 ( .A(msg[27]), .Y(n13719) );
  INVX1 U8216 ( .A(msg[30]), .Y(n13708) );
  AOI22X1 U8217 ( .A(msg[30]), .B(n13719), .C(msg[27]), .D(n13708), .Y(n13308)
         );
  XNOR2X1 U8218 ( .A(n11398), .B(n11150), .Y(n11605) );
  INVX1 U8219 ( .A(msg[2]), .Y(n13811) );
  INVX1 U8220 ( .A(msg[5]), .Y(n13799) );
  INVX1 U8221 ( .A(msg[33]), .Y(n13683) );
  MUX2X1 U8222 ( .B(msg[5]), .A(n13799), .S(n13683), .Y(n11393) );
  MUX2X1 U8223 ( .B(msg[2]), .A(n13811), .S(n11393), .Y(n12640) );
  XNOR2X1 U8224 ( .A(n11241), .B(n12640), .Y(n11576) );
  INVX1 U8225 ( .A(msg[13]), .Y(n13764) );
  MUX2X1 U8226 ( .B(msg[13]), .A(n13764), .S(n13775), .Y(n11388) );
  MUX2X1 U8227 ( .B(msg[25]), .A(n13723), .S(n11388), .Y(n11242) );
  FAX1 U8228 ( .A(msg[19]), .B(n11364), .C(n11242), .YS(n11243) );
  FAX1 U8229 ( .A(n11605), .B(n11576), .C(n11243), .YS(n11244) );
  FAX1 U8230 ( .A(n11319), .B(n11339), .C(n11244), .YS(n11474) );
  OR2X1 U8231 ( .A(n11474), .B(n11712), .Y(n12675) );
  AND2X1 U8232 ( .A(n10689), .B(n12675), .Y(n12677) );
  INVX1 U8233 ( .A(msg[53]), .Y(n11245) );
  AOI22X1 U8234 ( .A(msg[53]), .B(n13711), .C(msg[29]), .D(n11245), .Y(n12652)
         );
  INVX1 U8235 ( .A(n11167), .Y(n12651) );
  HAX1 U8236 ( .A(n12651), .B(n11591), .YS(n11246) );
  FAX1 U8237 ( .A(n11247), .B(n11388), .C(n11246), .YS(n11400) );
  INVX1 U8238 ( .A(msg[50]), .Y(n11273) );
  INVX1 U8239 ( .A(msg[41]), .Y(n13646) );
  MUX2X1 U8240 ( .B(msg[41]), .A(n13646), .S(n13731), .Y(n11281) );
  MUX2X1 U8241 ( .B(n11273), .A(msg[50]), .S(n11281), .Y(n11593) );
  MUX2X1 U8242 ( .B(n13783), .A(msg[9]), .S(n11593), .Y(n11372) );
  AOI22X1 U8243 ( .A(msg[32]), .B(msg[15]), .C(n13758), .D(n13688), .Y(n11248)
         );
  FAX1 U8244 ( .A(n11249), .B(n11191), .C(n10692), .YS(n11253) );
  INVX1 U8245 ( .A(msg[35]), .Y(n13679) );
  INVX1 U8246 ( .A(msg[47]), .Y(n11285) );
  INVX1 U8247 ( .A(msg[38]), .Y(n13671) );
  MUX2X1 U8248 ( .B(msg[18]), .A(n13737), .S(n13671), .Y(n11258) );
  MUX2X1 U8249 ( .B(n11285), .A(msg[47]), .S(n11258), .Y(n12638) );
  INVX1 U8250 ( .A(n12638), .Y(n12639) );
  HAX1 U8251 ( .A(n13299), .B(n12639), .YS(n11347) );
  INVX1 U8252 ( .A(msg[56]), .Y(n11351) );
  MUX2X1 U8253 ( .B(msg[24]), .A(n13725), .S(n11351), .Y(n11250) );
  FAX1 U8254 ( .A(msg[44]), .B(n11347), .C(n11250), .YS(n11251) );
  MUX2X1 U8255 ( .B(msg[35]), .A(n13679), .S(n11251), .Y(n11252) );
  FAX1 U8256 ( .A(n11254), .B(n11253), .C(n11252), .YS(n11255) );
  FAX1 U8257 ( .A(n11400), .B(n11372), .C(n11255), .YS(n11711) );
  INVX1 U8258 ( .A(msg[57]), .Y(n11338) );
  MUX2X1 U8259 ( .B(msg[57]), .A(n11338), .S(n12641), .Y(n11280) );
  MUX2X1 U8260 ( .B(n13729), .A(msg[22]), .S(n11281), .Y(n12649) );
  INVX1 U8261 ( .A(msg[44]), .Y(n11267) );
  MUX2X1 U8262 ( .B(n11267), .A(msg[44]), .S(n13625), .Y(n11590) );
  XNOR2X1 U8263 ( .A(n11388), .B(n11590), .Y(n11366) );
  MUX2X1 U8264 ( .B(msg[20]), .A(n13733), .S(n13761), .Y(n11256) );
  MUX2X1 U8265 ( .B(n13683), .A(msg[33]), .S(n11256), .Y(n11257) );
  MUX2X1 U8266 ( .B(n13677), .A(msg[36]), .S(n11257), .Y(n11264) );
  INVX1 U8267 ( .A(msg[54]), .Y(n11595) );
  MUX2X1 U8268 ( .B(n11595), .A(msg[54]), .S(n11258), .Y(n11278) );
  INVX1 U8269 ( .A(msg[51]), .Y(n11571) );
  MUX2X1 U8270 ( .B(msg[35]), .A(n13679), .S(n11096), .Y(n11348) );
  MUX2X1 U8271 ( .B(n11571), .A(msg[51]), .S(n11348), .Y(n11316) );
  INVX1 U8272 ( .A(msg[0]), .Y(n13821) );
  MUX2X1 U8273 ( .B(n13821), .A(msg[0]), .S(n11288), .Y(n11588) );
  HAX1 U8274 ( .A(n11316), .B(n11588), .YS(n11260) );
  MUX2X1 U8275 ( .B(n13725), .A(msg[24]), .S(n11260), .Y(n11375) );
  MUX2X1 U8276 ( .B(n13739), .A(msg[17]), .S(n11605), .Y(n11261) );
  MUX2X1 U8277 ( .B(msg[16]), .A(n13743), .S(n11261), .Y(n11262) );
  FAX1 U8278 ( .A(n11278), .B(n11375), .C(n11262), .YS(n11263) );
  FAX1 U8279 ( .A(n11366), .B(n11264), .C(n11263), .YS(n11265) );
  FAX1 U8280 ( .A(n11280), .B(n12649), .C(n11265), .YS(n11709) );
  INVX1 U8281 ( .A(n11474), .Y(n13253) );
  NAND2X1 U8282 ( .A(n11010), .B(n13253), .Y(n11292) );
  OAI21X1 U8283 ( .A(n12677), .B(n11711), .C(n11292), .Y(n10379) );
  HAX1 U8284 ( .A(n11266), .B(n13306), .YS(n11318) );
  AOI22X1 U8285 ( .A(msg[52]), .B(msg[0]), .C(n13821), .D(n11336), .Y(n11268)
         );
  MUX2X1 U8286 ( .B(n12646), .A(msg[48]), .S(n11267), .Y(n11606) );
  FAX1 U8287 ( .A(n11094), .B(msg[56]), .C(n11606), .YS(n11269) );
  FAX1 U8288 ( .A(n11270), .B(n11318), .C(n11269), .YS(n13083) );
  MUX2X1 U8289 ( .B(n13708), .A(msg[30]), .S(n11271), .Y(n11272) );
  MUX2X1 U8290 ( .B(n13779), .A(msg[10]), .S(n11272), .Y(n11320) );
  INVX1 U8291 ( .A(n12645), .Y(n12644) );
  MUX2X1 U8292 ( .B(msg[26]), .A(n13721), .S(n11273), .Y(n11274) );
  MUX2X1 U8293 ( .B(n13795), .A(msg[6]), .S(n11274), .Y(n11275) );
  MUX2X1 U8294 ( .B(msg[2]), .A(n13811), .S(n11275), .Y(n11276) );
  FAX1 U8295 ( .A(n12644), .B(n11384), .C(n11276), .YS(n11277) );
  FAX1 U8296 ( .A(n11278), .B(n11320), .C(n11277), .YS(n12685) );
  NAND2X1 U8297 ( .A(n13083), .B(n12685), .Y(n11394) );
  HAX1 U8298 ( .A(n11280), .B(n11279), .YS(n11574) );
  MUX2X1 U8299 ( .B(n13764), .A(msg[13]), .S(n11393), .Y(n11613) );
  MUX2X1 U8300 ( .B(n13815), .A(msg[1]), .S(n11281), .Y(n11282) );
  FAX1 U8301 ( .A(n11282), .B(n11369), .C(n11167), .YS(n11283) );
  FAX1 U8302 ( .A(n11574), .B(n11613), .C(n11283), .YS(n13085) );
  MUX2X1 U8303 ( .B(n11285), .A(msg[47]), .S(n11284), .Y(n11286) );
  MUX2X1 U8304 ( .B(n13807), .A(msg[3]), .S(n11286), .Y(n11287) );
  MUX2X1 U8305 ( .B(n13705), .A(msg[31]), .S(n11287), .Y(n11627) );
  MUX2X1 U8306 ( .B(n13679), .A(msg[35]), .S(n11288), .Y(n11343) );
  MUX2X1 U8307 ( .B(msg[27]), .A(n13719), .S(n13300), .Y(n11289) );
  MUX2X1 U8308 ( .B(n13791), .A(msg[7]), .S(n11289), .Y(n12637) );
  AOI22X1 U8309 ( .A(msg[15]), .B(n13727), .C(msg[23]), .D(n13758), .Y(n11290)
         );
  FAX1 U8310 ( .A(n12637), .B(msg[51]), .C(n10693), .YS(n11291) );
  FAX1 U8311 ( .A(n11627), .B(n11343), .C(n11291), .YS(n12696) );
  AND2X1 U8312 ( .A(n12682), .B(n10379), .Y(
        \lamb/scale_ts1/genblk1[3].mult/logA[0] ) );
  AND2X1 U8313 ( .A(n11712), .B(n11711), .Y(n11293) );
  AOI22X1 U8314 ( .A(n11010), .B(n11474), .C(n11712), .D(n11711), .Y(n11294)
         );
  INVX1 U8315 ( .A(n11711), .Y(n12679) );
  OAI21X1 U8316 ( .A(n13255), .B(n11294), .C(n13259), .Y(
        \lamb/scale_ts0/genblk1[2].mult/logA[2] ) );
  AND2X1 U8317 ( .A(n12682), .B(\lamb/scale_ts0/genblk1[2].mult/logA[2] ), .Y(
        \lamb/scale_ls2/genblk1[1].mult/logA[2] ) );
  INVX1 U8318 ( .A(\lamb/scale_ds1/genblk1[3].mult/added[4] ), .Y(n11296) );
  NAND2X1 U8319 ( .A(\add_x_146/n1 ), .B(
        \lamb/scale_ds1/genblk1[3].mult/added[3] ), .Y(n11302) );
  INVX1 U8320 ( .A(\lamb/scale_ds1/genblk1[3].mult/added[3] ), .Y(n11297) );
  NAND2X1 U8321 ( .A(n11297), .B(n11296), .Y(n11304) );
  INVX1 U8322 ( .A(\lamb/scale_ds1/genblk1[3].mult/added[2] ), .Y(n11427) );
  INVX1 U8323 ( .A(\lamb/scale_ds1/genblk1[3].mult/added[1] ), .Y(n11298) );
  NOR2X1 U8324 ( .A(n11427), .B(n11298), .Y(n11295) );
  OAI21X1 U8325 ( .A(n10668), .B(n11295), .C(n11300), .Y(n11456) );
  OAI21X1 U8326 ( .A(\lamb/scale_ds1/genblk1[3].mult/added[1] ), .B(n10423), 
        .C(n11456), .Y(n11383) );
  OR2X1 U8327 ( .A(n11427), .B(n10668), .Y(n11429) );
  INVX1 U8328 ( .A(n11429), .Y(n11307) );
  INVX1 U8329 ( .A(\add_x_146/n1 ), .Y(n11301) );
  AOI22X1 U8330 ( .A(\add_x_146/n1 ), .B(n11296), .C(
        \lamb/scale_ds1/genblk1[3].mult/added[4] ), .D(n11301), .Y(n11430) );
  NOR2X1 U8331 ( .A(n11297), .B(n11430), .Y(n11299) );
  NOR2X1 U8332 ( .A(\lamb/scale_ds1/genblk1[3].mult/added[2] ), .B(n11106), 
        .Y(n11306) );
  NAND3X1 U8333 ( .A(n11304), .B(n10940), .C(n11302), .Y(n11425) );
  INVX1 U8334 ( .A(n11425), .Y(n11437) );
  NAND2X1 U8335 ( .A(\lamb/scale_ds1/genblk1[3].mult/added[1] ), .B(n11437), 
        .Y(n11305) );
  AOI22X1 U8336 ( .A(n11307), .B(n11052), .C(n11306), .D(n11305), .Y(n11461)
         );
  INVX1 U8337 ( .A(\lamb/scale_ts0/genblk1[2].mult/added[1] ), .Y(n11379) );
  NAND2X1 U8338 ( .A(\lamb/scale_ts0/genblk1[2].mult/added[2] ), .B(n11379), 
        .Y(n11309) );
  NAND3X1 U8339 ( .A(\lamb/scale_ts0/genblk1[2].mult/added[3] ), .B(n10669), 
        .C(n11329), .Y(n11323) );
  INVX1 U8340 ( .A(\lamb/scale_ts0/genblk1[2].mult/added[3] ), .Y(n11327) );
  INVX1 U8341 ( .A(\lamb/scale_ts0/genblk1[2].mult/added[2] ), .Y(n11330) );
  AOI22X1 U8342 ( .A(\lamb/scale_ts0/genblk1[2].mult/added[2] ), .B(n11308), 
        .C(n11123), .D(n11330), .Y(n11325) );
  OAI21X1 U8343 ( .A(n11309), .B(n11323), .C(n11325), .Y(n11381) );
  NAND3X1 U8344 ( .A(n11123), .B(\lamb/scale_ts0/genblk1[2].mult/added[2] ), 
        .C(n11379), .Y(n11334) );
  NOR2X1 U8345 ( .A(n11379), .B(n11330), .Y(n11311) );
  AOI22X1 U8346 ( .A(n11311), .B(n11310), .C(n11173), .D(n11327), .Y(n11376)
         );
  NAND3X1 U8347 ( .A(\lamb/scale_ts0/genblk1[2].mult/added[4] ), .B(
        \add_x_152/n1 ), .C(n11327), .Y(n11312) );
  OAI21X1 U8348 ( .A(n11329), .B(n11327), .C(n11312), .Y(n11328) );
  NAND2X1 U8349 ( .A(\lamb/scale_ts0/genblk1[2].mult/added[1] ), .B(n11328), 
        .Y(n11313) );
  NAND3X1 U8350 ( .A(n11334), .B(n11376), .C(n11313), .Y(n11315) );
  NAND2X1 U8351 ( .A(n10689), .B(n11711), .Y(n12674) );
  INVX1 U8352 ( .A(n12674), .Y(n11314) );
  NOR2X1 U8353 ( .A(n11010), .B(n13253), .Y(n12680) );
  OAI21X1 U8354 ( .A(n11381), .B(n11315), .C(n11857), .Y(n11322) );
  MUX2X1 U8355 ( .B(msg[1]), .A(n13815), .S(n11316), .Y(n11317) );
  XNOR2X1 U8356 ( .A(n11318), .B(n11317), .Y(n11633) );
  HAX1 U8357 ( .A(n11320), .B(n11319), .YS(n11598) );
  MUX2X1 U8358 ( .B(msg[41]), .A(n13646), .S(msg[53]), .Y(n11390) );
  MUX2X1 U8359 ( .B(msg[39]), .A(n13669), .S(n11390), .Y(n13303) );
  FAX1 U8360 ( .A(msg[45]), .B(n11576), .C(n13303), .YS(n11321) );
  FAX1 U8361 ( .A(n11633), .B(n11598), .C(n11321), .YS(n12293) );
  INVX1 U8362 ( .A(n12293), .Y(n13372) );
  HAX1 U8363 ( .A(n11322), .B(n13372), .YS(n13834) );
  INVX1 U8364 ( .A(n13834), .Y(n13332) );
  NAND2X1 U8365 ( .A(\lamb/scale_ts0/genblk1[2].mult/added[2] ), .B(n11328), 
        .Y(n11360) );
  NAND2X1 U8366 ( .A(n11379), .B(n11360), .Y(n11333) );
  INVX1 U8367 ( .A(n11323), .Y(n11359) );
  NAND3X1 U8368 ( .A(\lamb/scale_ts0/genblk1[2].mult/added[1] ), .B(n11325), 
        .C(n10964), .Y(n11356) );
  NAND3X1 U8369 ( .A(n11327), .B(n10669), .C(n11329), .Y(n11378) );
  AOI21X1 U8370 ( .A(\lamb/scale_ts0/genblk1[2].mult/added[1] ), .B(n11173), 
        .C(n11328), .Y(n11331) );
  AOI22X1 U8371 ( .A(\lamb/scale_ts0/genblk1[2].mult/added[2] ), .B(n10656), 
        .C(n11331), .D(n11330), .Y(n11332) );
  AOI21X1 U8372 ( .A(n11333), .B(n11356), .C(n11332), .Y(n11335) );
  AOI21X1 U8373 ( .A(n11335), .B(n11334), .C(n10799), .Y(n11346) );
  MUX2X1 U8374 ( .B(n11336), .A(msg[52]), .S(n11593), .Y(n11397) );
  MUX2X1 U8375 ( .B(msg[5]), .A(n13799), .S(n11397), .Y(n11631) );
  INVX1 U8376 ( .A(n11631), .Y(n11345) );
  HAX1 U8377 ( .A(n12639), .B(n11337), .YS(n11615) );
  MUX2X1 U8378 ( .B(msg[57]), .A(n11338), .S(msg[55]), .Y(n13296) );
  MUX2X1 U8379 ( .B(msg[37]), .A(n13673), .S(n13296), .Y(n11342) );
  FAX1 U8380 ( .A(msg[45]), .B(n11398), .C(n11339), .YS(n11340) );
  MUX2X1 U8381 ( .B(msg[26]), .A(n13721), .S(n11340), .Y(n11341) );
  FAX1 U8382 ( .A(n11343), .B(n11342), .C(n11341), .YS(n11344) );
  FAX1 U8383 ( .A(n11345), .B(n11615), .C(n11344), .YS(n11568) );
  INVX1 U8384 ( .A(n11568), .Y(n13370) );
  HAX1 U8385 ( .A(n11346), .B(n13370), .YS(n13337) );
  INVX1 U8386 ( .A(n13337), .Y(n13837) );
  AND2X1 U8387 ( .A(n13332), .B(n13837), .Y(n13334) );
  FAX1 U8388 ( .A(n11160), .B(n11348), .C(n11347), .YS(n11350) );
  MUX2X1 U8389 ( .B(n13803), .A(msg[4]), .S(n11350), .Y(n11401) );
  AOI22X1 U8390 ( .A(msg[56]), .B(msg[23]), .C(n13727), .D(n11351), .Y(n11626)
         );
  MUX2X1 U8391 ( .B(n11595), .A(msg[54]), .S(msg[46]), .Y(n11608) );
  AOI22X1 U8392 ( .A(msg[34]), .B(msg[7]), .C(n13791), .D(n13681), .Y(n11352)
         );
  FAX1 U8393 ( .A(n11156), .B(n11608), .C(n10694), .YS(n11353) );
  MUX2X1 U8394 ( .B(msg[25]), .A(n13723), .S(n11353), .Y(n11354) );
  FAX1 U8395 ( .A(n11366), .B(n11587), .C(n11354), .YS(n11355) );
  FAX1 U8396 ( .A(n11401), .B(n11576), .C(n11355), .YS(n13826) );
  INVX1 U8397 ( .A(n13826), .Y(n13377) );
  INVX1 U8398 ( .A(n11356), .Y(n11357) );
  NAND2X1 U8399 ( .A(n11357), .B(n10656), .Y(n11358) );
  OAI21X1 U8400 ( .A(\lamb/scale_ts0/genblk1[2].mult/added[1] ), .B(n11359), 
        .C(n11358), .Y(n11361) );
  NAND2X1 U8401 ( .A(n10898), .B(n11857), .Y(n11363) );
  HAX1 U8402 ( .A(n13377), .B(n11363), .YS(n13830) );
  MUX2X1 U8403 ( .B(n13719), .A(msg[27]), .S(n11364), .Y(n11365) );
  MUX2X1 U8404 ( .B(n13795), .A(msg[6]), .S(n11365), .Y(n11374) );
  HAX1 U8405 ( .A(n12651), .B(n11366), .YS(n11367) );
  MUX2X1 U8406 ( .B(n13770), .A(msg[12]), .S(n11367), .Y(n11573) );
  MUX2X1 U8407 ( .B(n13787), .A(msg[8]), .S(msg[58]), .Y(n11607) );
  HAX1 U8408 ( .A(n11369), .B(n11191), .YS(n13302) );
  FAX1 U8409 ( .A(msg[38]), .B(n11607), .C(n13302), .YS(n11370) );
  MUX2X1 U8410 ( .B(msg[40]), .A(n13666), .S(n11370), .Y(n11371) );
  FAX1 U8411 ( .A(n11372), .B(n11573), .C(n11371), .YS(n11373) );
  FAX1 U8412 ( .A(n11375), .B(n11374), .C(n11373), .YS(n13367) );
  INVX1 U8413 ( .A(n13367), .Y(n13371) );
  INVX1 U8414 ( .A(n11376), .Y(n11377) );
  AOI21X1 U8415 ( .A(n11379), .B(n10656), .C(n11377), .Y(n11380) );
  OAI21X1 U8416 ( .A(n11381), .B(n10939), .C(n11857), .Y(n11382) );
  HAX1 U8417 ( .A(n13371), .B(n11382), .YS(n13336) );
  NAND3X1 U8418 ( .A(n13334), .B(n13830), .C(n13336), .Y(n11459) );
  OAI21X1 U8419 ( .A(n11383), .B(n10385), .C(n11152), .Y(n11410) );
  MUX2X1 U8420 ( .B(n13705), .A(msg[31]), .S(n11384), .Y(n11385) );
  MUX2X1 U8421 ( .B(msg[9]), .A(n13783), .S(n11385), .Y(n11386) );
  FAX1 U8422 ( .A(msg[57]), .B(n11387), .C(n11386), .YS(n11389) );
  FAX1 U8423 ( .A(n11390), .B(n11389), .C(n11388), .YS(n11391) );
  FAX1 U8424 ( .A(n11393), .B(n11392), .C(n11391), .YS(n13325) );
  INVX1 U8425 ( .A(n13083), .Y(n13225) );
  INVX1 U8426 ( .A(n12685), .Y(n13231) );
  AOI22X1 U8427 ( .A(msg[0]), .B(n13783), .C(msg[9]), .D(n13821), .Y(n11396)
         );
  FAX1 U8428 ( .A(n11398), .B(n11397), .C(n10695), .YS(n11399) );
  FAX1 U8429 ( .A(n11401), .B(n11400), .C(n11399), .YS(n13317) );
  INVX1 U8430 ( .A(n13224), .Y(n12695) );
  INVX1 U8431 ( .A(n13085), .Y(n13229) );
  INVX1 U8432 ( .A(n12696), .Y(n12760) );
  HAX1 U8433 ( .A(n13253), .B(n10674), .YS(n13324) );
  NAND2X1 U8434 ( .A(n12695), .B(n13324), .Y(n12304) );
  AND2X1 U8435 ( .A(\add_x_142/n1 ), .B(
        \lamb/scale_ts1/genblk1[3].mult/added[4] ), .Y(n11404) );
  OR2X1 U8436 ( .A(n10672), .B(\lamb/scale_ts1/genblk1[3].mult/added[1] ), .Y(
        n11420) );
  NAND2X1 U8437 ( .A(\lamb/scale_ts1/genblk1[3].mult/added[1] ), .B(
        \lamb/scale_ts1/genblk1[3].mult/added[2] ), .Y(n11414) );
  INVX1 U8438 ( .A(n11414), .Y(n11402) );
  OR2X1 U8439 ( .A(\add_x_142/n1 ), .B(
        \lamb/scale_ts1/genblk1[3].mult/added[4] ), .Y(n11419) );
  AOI21X1 U8440 ( .A(n11402), .B(n10672), .C(n10666), .Y(n11451) );
  AOI21X1 U8441 ( .A(\add_x_142/n1 ), .B(
        \lamb/scale_ts1/genblk1[3].mult/added[4] ), .C(
        \lamb/scale_ts1/genblk1[3].mult/added[3] ), .Y(n11452) );
  INVX1 U8442 ( .A(n10552), .Y(n11411) );
  NOR3X1 U8443 ( .A(\lamb/scale_ts1/genblk1[3].mult/added[1] ), .B(n11404), 
        .C(n10734), .Y(n11442) );
  OAI21X1 U8444 ( .A(n10666), .B(n11442), .C(
        \lamb/scale_ts1/genblk1[3].mult/added[2] ), .Y(n11405) );
  OAI21X1 U8445 ( .A(\lamb/scale_ts1/genblk1[3].mult/added[2] ), .B(n10672), 
        .C(n11405), .Y(n11415) );
  INVX1 U8446 ( .A(n11415), .Y(n11455) );
  NAND3X1 U8447 ( .A(n11420), .B(n11407), .C(n11455), .Y(n11408) );
  NAND2X1 U8448 ( .A(n11453), .B(n11408), .Y(n11409) );
  HAX1 U8449 ( .A(n11410), .B(n11409), .YS(n13846) );
  INVX1 U8450 ( .A(n13846), .Y(n13854) );
  NAND2X1 U8451 ( .A(\lamb/scale_ts1/genblk1[3].mult/added[2] ), .B(n11416), 
        .Y(n11443) );
  OAI21X1 U8452 ( .A(n10734), .B(n10902), .C(n11443), .Y(n11413) );
  AOI22X1 U8453 ( .A(\lamb/scale_ts1/genblk1[3].mult/added[1] ), .B(n11415), 
        .C(n11414), .D(n11413), .Y(n11447) );
  AOI21X1 U8454 ( .A(n10666), .B(\lamb/scale_ts1/genblk1[3].mult/added[1] ), 
        .C(n11416), .Y(n11418) );
  INVX1 U8455 ( .A(n11418), .Y(n11422) );
  NAND3X1 U8456 ( .A(n11050), .B(n11420), .C(
        \lamb/scale_ts1/genblk1[3].mult/added[2] ), .Y(n11421) );
  OAI21X1 U8457 ( .A(\lamb/scale_ts1/genblk1[3].mult/added[2] ), .B(n11422), 
        .C(n11421), .Y(n11423) );
  AOI21X1 U8458 ( .A(n11447), .B(n11423), .C(n11115), .Y(n11436) );
  AOI22X1 U8459 ( .A(\lamb/scale_ds1/genblk1[3].mult/added[2] ), .B(
        \lamb/scale_ds1/genblk1[3].mult/added[1] ), .C(n11425), .D(n10423), 
        .Y(n11434) );
  OAI21X1 U8460 ( .A(\lamb/scale_ds1/genblk1[3].mult/added[4] ), .B(
        \add_x_146/n1 ), .C(\lamb/scale_ds1/genblk1[3].mult/added[3] ), .Y(
        n11426) );
  NAND3X1 U8461 ( .A(\lamb/scale_ds1/genblk1[3].mult/added[1] ), .B(n11429), 
        .C(n10958), .Y(n11438) );
  AOI22X1 U8462 ( .A(n10668), .B(\lamb/scale_ds1/genblk1[3].mult/added[1] ), 
        .C(\lamb/scale_ds1/genblk1[3].mult/added[2] ), .D(n11144), .Y(n11432)
         );
  NAND2X1 U8463 ( .A(n11438), .B(n11432), .Y(n11433) );
  OAI21X1 U8464 ( .A(n11434), .B(n11433), .C(n11152), .Y(n11435) );
  HAX1 U8465 ( .A(n11436), .B(n11435), .YS(n13855) );
  AOI22X1 U8466 ( .A(\lamb/scale_ds1/genblk1[3].mult/added[2] ), .B(n11437), 
        .C(\lamb/scale_ds1/genblk1[3].mult/added[1] ), .D(n11144), .Y(n11439)
         );
  NAND3X1 U8467 ( .A(n11052), .B(n11439), .C(n11438), .Y(n11441) );
  NAND2X1 U8468 ( .A(n11441), .B(n11152), .Y(n11450) );
  AOI21X1 U8469 ( .A(n11050), .B(n11443), .C(n10902), .Y(n11445) );
  INVX1 U8470 ( .A(n11445), .Y(n11446) );
  NAND2X1 U8471 ( .A(n11453), .B(n11448), .Y(n11449) );
  HAX1 U8472 ( .A(n11450), .B(n11449), .YS(n13857) );
  INVX1 U8473 ( .A(n13857), .Y(n13852) );
  AND2X1 U8474 ( .A(n13855), .B(n13852), .Y(n13840) );
  OAI21X1 U8475 ( .A(\lamb/scale_ts1/genblk1[3].mult/added[1] ), .B(n10552), 
        .C(n10994), .Y(n11454) );
  AOI21X1 U8476 ( .A(n11455), .B(n11454), .C(n11115), .Y(n11464) );
  OAI21X1 U8477 ( .A(\lamb/scale_ds1/genblk1[3].mult/added[1] ), .B(n11144), 
        .C(n11456), .Y(n11458) );
  INVX1 U8478 ( .A(n11458), .Y(n11460) );
  OAI21X1 U8479 ( .A(n10385), .B(n11460), .C(n11152), .Y(n11462) );
  INVX1 U8480 ( .A(n11462), .Y(n11463) );
  HAX1 U8481 ( .A(n11464), .B(n11463), .YS(n13850) );
  INVX1 U8482 ( .A(n13850), .Y(n13848) );
  INVX1 U8483 ( .A(n10591), .Y(n12698) );
  NAND2X1 U8484 ( .A(n13854), .B(n12698), .Y(n12215) );
  NAND2X1 U8485 ( .A(n12682), .B(n12215), .Y(n11511) );
  INVX1 U8486 ( .A(n11511), .Y(n11534) );
  AOI21X1 U8487 ( .A(\lamb/scale_bs2/genblk1[0].mult/added[4] ), .B(
        \add_x_138/n1 ), .C(n10825), .Y(n11517) );
  AND2X1 U8488 ( .A(\lamb/scale_bs2/genblk1[0].mult/added[2] ), .B(n10815), 
        .Y(n11468) );
  INVX1 U8489 ( .A(\lamb/scale_bs2/genblk1[0].mult/added[3] ), .Y(n11514) );
  NAND2X1 U8490 ( .A(\lamb/scale_bs2/genblk1[0].mult/added[2] ), .B(
        \lamb/scale_bs2/genblk1[0].mult/added[1] ), .Y(n11515) );
  AND2X1 U8491 ( .A(\add_x_138/n1 ), .B(
        \lamb/scale_bs2/genblk1[0].mult/added[4] ), .Y(n11465) );
  AOI22X1 U8492 ( .A(\lamb/scale_bs2/genblk1[0].mult/added[3] ), .B(n10825), 
        .C(n11465), .D(n11514), .Y(n11518) );
  NAND3X1 U8493 ( .A(\lamb/scale_bs2/genblk1[0].mult/added[2] ), .B(n11465), 
        .C(\lamb/scale_bs2/genblk1[0].mult/added[3] ), .Y(n11499) );
  OAI21X1 U8494 ( .A(n10825), .B(\lamb/scale_bs2/genblk1[0].mult/added[3] ), 
        .C(\lamb/scale_bs2/genblk1[0].mult/added[1] ), .Y(n11466) );
  NAND3X1 U8495 ( .A(n11107), .B(n10700), .C(n11466), .Y(n11467) );
  AOI22X1 U8496 ( .A(n11468), .B(n11514), .C(n11515), .D(n11467), .Y(n11473)
         );
  INVX1 U8497 ( .A(\lamb/scale_bs2/genblk1[0].mult/added[1] ), .Y(n11519) );
  NAND3X1 U8498 ( .A(\lamb/scale_bs2/genblk1[0].mult/added[3] ), .B(n10815), 
        .C(n11519), .Y(n11470) );
  NAND2X1 U8499 ( .A(n10825), .B(n11514), .Y(n11469) );
  NAND3X1 U8500 ( .A(\lamb/scale_bs2/genblk1[0].mult/added[2] ), .B(n11470), 
        .C(n11469), .Y(n11503) );
  INVX1 U8501 ( .A(\lamb/scale_bs2/genblk1[0].mult/added[2] ), .Y(n11472) );
  NAND3X1 U8502 ( .A(\add_x_138/n1 ), .B(
        \lamb/scale_bs2/genblk1[0].mult/added[4] ), .C(
        \lamb/scale_bs2/genblk1[0].mult/added[3] ), .Y(n11471) );
  NAND2X1 U8503 ( .A(n11472), .B(n11471), .Y(n11484) );
  NAND2X1 U8504 ( .A(n11474), .B(n12695), .Y(n11714) );
  NOR2X1 U8505 ( .A(\add_x_141/n1 ), .B(
        \lamb/scale_ls2/genblk1[0].mult/added[4] ), .Y(n11476) );
  AOI21X1 U8506 ( .A(\lamb/scale_ls2/genblk1[0].mult/added[4] ), .B(
        \add_x_141/n1 ), .C(n11476), .Y(n11505) );
  INVX1 U8507 ( .A(\lamb/scale_ls2/genblk1[0].mult/added[3] ), .Y(n11475) );
  INVX1 U8508 ( .A(\lamb/scale_ls2/genblk1[0].mult/added[1] ), .Y(n11494) );
  AND2X1 U8509 ( .A(\lamb/scale_ls2/genblk1[0].mult/added[2] ), .B(n10621), 
        .Y(n11528) );
  OAI21X1 U8510 ( .A(n11494), .B(n11528), .C(n10660), .Y(n11477) );
  OAI21X1 U8511 ( .A(\lamb/scale_ls2/genblk1[0].mult/added[2] ), .B(n10660), 
        .C(n11477), .Y(n11481) );
  AND2X1 U8512 ( .A(\add_x_141/n1 ), .B(
        \lamb/scale_ls2/genblk1[0].mult/added[4] ), .Y(n11478) );
  NAND3X1 U8513 ( .A(\lamb/scale_ls2/genblk1[0].mult/added[2] ), .B(n11526), 
        .C(n11494), .Y(n11507) );
  NOR2X1 U8514 ( .A(n11159), .B(n11526), .Y(n11479) );
  NAND3X1 U8515 ( .A(n11479), .B(n11494), .C(n10621), .Y(n11480) );
  NAND3X1 U8516 ( .A(n11481), .B(n11085), .C(n11480), .Y(n11482) );
  AOI22X1 U8517 ( .A(n11534), .B(n10927), .C(n13258), .D(n11482), .Y(n11513)
         );
  AOI21X1 U8518 ( .A(n10825), .B(n11514), .C(n11484), .Y(n11486) );
  INVX1 U8519 ( .A(n11486), .Y(n11502) );
  AOI21X1 U8520 ( .A(n10700), .B(n11502), .C(n11519), .Y(n11487) );
  INVX1 U8521 ( .A(n11487), .Y(n11490) );
  NAND3X1 U8522 ( .A(n10815), .B(n11514), .C(n11519), .Y(n11488) );
  NAND3X1 U8523 ( .A(n11490), .B(n11048), .C(n11488), .Y(n11497) );
  NAND3X1 U8524 ( .A(n11159), .B(\lamb/scale_ls2/genblk1[0].mult/added[3] ), 
        .C(n11494), .Y(n11531) );
  INVX1 U8525 ( .A(\lamb/scale_ls2/genblk1[0].mult/added[2] ), .Y(n11506) );
  AOI22X1 U8526 ( .A(n11528), .B(n11531), .C(n11506), .D(n10783), .Y(n11525)
         );
  NAND3X1 U8527 ( .A(\lamb/scale_ls2/genblk1[0].mult/added[2] ), .B(
        \lamb/scale_ls2/genblk1[0].mult/added[1] ), .C(n10783), .Y(n11491) );
  AOI21X1 U8528 ( .A(n11494), .B(n10660), .C(n10990), .Y(n11495) );
  OR2X1 U8529 ( .A(n10670), .B(n11495), .Y(n11496) );
  AOI22X1 U8530 ( .A(n11534), .B(n11497), .C(n13258), .D(n11496), .Y(n13137)
         );
  INVX1 U8531 ( .A(n11107), .Y(n11498) );
  AOI21X1 U8532 ( .A(\lamb/scale_bs2/genblk1[0].mult/added[2] ), .B(n10815), 
        .C(n11498), .Y(n11500) );
  AOI22X1 U8533 ( .A(\lamb/scale_bs2/genblk1[0].mult/added[1] ), .B(n11500), 
        .C(n10700), .D(n11519), .Y(n11501) );
  AOI21X1 U8534 ( .A(n11503), .B(n11502), .C(n10909), .Y(n11512) );
  INVX1 U8535 ( .A(n11159), .Y(n11527) );
  NAND3X1 U8536 ( .A(\lamb/scale_ls2/genblk1[0].mult/added[1] ), .B(n11527), 
        .C(n11506), .Y(n11508) );
  NAND3X1 U8537 ( .A(n11504), .B(n11508), .C(n11085), .Y(n11509) );
  OAI21X1 U8538 ( .A(n10670), .B(n11509), .C(n13258), .Y(n11510) );
  OAI21X1 U8539 ( .A(n11512), .B(n11511), .C(n11510), .Y(n12767) );
  NAND2X1 U8540 ( .A(n10483), .B(n12767), .Y(n12768) );
  AND2X1 U8541 ( .A(n11513), .B(n12768), .Y(n13147) );
  INVX1 U8542 ( .A(n10483), .Y(n13141) );
  INVX1 U8543 ( .A(n11513), .Y(n13143) );
  NAND2X1 U8544 ( .A(n11514), .B(n11519), .Y(n11516) );
  OAI21X1 U8545 ( .A(n11519), .B(\lamb/scale_bs2/genblk1[0].mult/added[3] ), 
        .C(n11107), .Y(n11520) );
  NAND2X1 U8546 ( .A(\lamb/scale_bs2/genblk1[0].mult/added[2] ), .B(n11520), 
        .Y(n11521) );
  NAND3X1 U8547 ( .A(n11523), .B(n11522), .C(n11521), .Y(n11533) );
  AOI21X1 U8548 ( .A(\lamb/scale_ls2/genblk1[0].mult/added[3] ), .B(
        \lamb/scale_ls2/genblk1[0].mult/added[2] ), .C(n11527), .Y(n11524) );
  OAI21X1 U8549 ( .A(n10670), .B(n11524), .C(
        \lamb/scale_ls2/genblk1[0].mult/added[1] ), .Y(n11530) );
  NAND3X1 U8550 ( .A(n11528), .B(n11527), .C(n10783), .Y(n11529) );
  NAND3X1 U8551 ( .A(n11531), .B(n11530), .C(n11529), .Y(n11532) );
  AOI22X1 U8552 ( .A(n11534), .B(n11533), .C(n13258), .D(n11532), .Y(n13150)
         );
  AOI21X1 U8553 ( .A(n13141), .B(n11177), .C(n10819), .Y(n13138) );
  NAND2X1 U8554 ( .A(\lamb/scale_ls3/genblk1[0].mult/added[1] ), .B(
        \lamb/scale_ls3/genblk1[0].mult/added[2] ), .Y(n11801) );
  INVX1 U8555 ( .A(n11801), .Y(n11535) );
  NAND2X1 U8556 ( .A(\lamb/scale_ls3/genblk1[0].mult/added[3] ), .B(n11542), 
        .Y(n11536) );
  OR2X1 U8557 ( .A(\add_x_128/n1 ), .B(
        \lamb/scale_ls3/genblk1[0].mult/added[4] ), .Y(n11543) );
  INVX1 U8558 ( .A(n11543), .Y(n11910) );
  INVX1 U8559 ( .A(\lamb/scale_ls3/genblk1[0].mult/added[3] ), .Y(n11541) );
  AOI22X1 U8560 ( .A(n11535), .B(n11536), .C(n11910), .D(n11541), .Y(n11802)
         );
  INVX1 U8561 ( .A(n11536), .Y(n11914) );
  NOR2X1 U8562 ( .A(n11541), .B(n11910), .Y(n11538) );
  INVX1 U8563 ( .A(\lamb/scale_ls3/genblk1[0].mult/added[1] ), .Y(n11537) );
  NAND3X1 U8564 ( .A(n11538), .B(n11537), .C(n11131), .Y(n11992) );
  NAND2X1 U8565 ( .A(n11910), .B(n11541), .Y(n11539) );
  NAND3X1 U8566 ( .A(n11992), .B(n11539), .C(
        \lamb/scale_ls3/genblk1[0].mult/added[2] ), .Y(n11540) );
  OAI21X1 U8567 ( .A(\lamb/scale_ls3/genblk1[0].mult/added[2] ), .B(n11914), 
        .C(n11540), .Y(n11804) );
  AOI22X1 U8568 ( .A(\lamb/scale_ls3/genblk1[0].mult/added[3] ), .B(n11543), 
        .C(n11131), .D(n11541), .Y(n11990) );
  INVX1 U8569 ( .A(n10588), .Y(n11915) );
  NAND2X1 U8570 ( .A(\lamb/scale_ls3/genblk1[0].mult/added[1] ), .B(n11915), 
        .Y(n11911) );
  OAI21X1 U8571 ( .A(\lamb/scale_ls3/genblk1[0].mult/added[1] ), .B(n11914), 
        .C(n11911), .Y(n11544) );
  NAND3X1 U8572 ( .A(n11051), .B(n11804), .C(n11544), .Y(n11545) );
  NAND2X1 U8573 ( .A(n10677), .B(n11545), .Y(n11794) );
  AOI21X1 U8574 ( .A(n10627), .B(n13846), .C(n10591), .Y(n13086) );
  INVX1 U8575 ( .A(n11227), .Y(n13841) );
  NAND2X1 U8576 ( .A(n10851), .B(n13253), .Y(n11646) );
  NOR3X1 U8577 ( .A(n10629), .B(\lamb/scale_ds2/genblk1[3].mult/added[3] ), 
        .C(n11759), .Y(n11773) );
  INVX1 U8578 ( .A(\lamb/scale_ds2/genblk1[3].mult/added[2] ), .Y(n11546) );
  INVX1 U8579 ( .A(\lamb/scale_ds2/genblk1[3].mult/added[3] ), .Y(n11760) );
  NOR2X1 U8580 ( .A(\lamb/scale_ds2/genblk1[3].mult/added[1] ), .B(n11548), 
        .Y(n11736) );
  NAND2X1 U8581 ( .A(n11736), .B(n11151), .Y(n11762) );
  NAND2X1 U8582 ( .A(n11760), .B(n11151), .Y(n11547) );
  NAND2X1 U8583 ( .A(n11548), .B(n11547), .Y(n11757) );
  NAND2X1 U8584 ( .A(n11762), .B(n11757), .Y(n11549) );
  AOI22X1 U8585 ( .A(n11773), .B(\lamb/scale_ds2/genblk1[3].mult/added[1] ), 
        .C(n11082), .D(n11549), .Y(n11707) );
  NAND2X1 U8586 ( .A(\lamb/scale_ds2/genblk1[3].mult/added[2] ), .B(n11168), 
        .Y(n11734) );
  NAND3X1 U8587 ( .A(\lamb/scale_ds2/genblk1[3].mult/added[1] ), .B(n11082), 
        .C(n11734), .Y(n11739) );
  OR2X1 U8588 ( .A(\lamb/scale_ds1/genblk1[2].mult/added[4] ), .B(
        \add_x_147/n1 ), .Y(n11676) );
  OR2X1 U8589 ( .A(n11676), .B(\lamb/scale_ds1/genblk1[2].mult/added[3] ), .Y(
        n11554) );
  NAND2X1 U8590 ( .A(\lamb/scale_ds1/genblk1[2].mult/added[2] ), .B(n11554), 
        .Y(n11672) );
  INVX1 U8591 ( .A(n11672), .Y(n11553) );
  NAND2X1 U8592 ( .A(\lamb/scale_ds1/genblk1[2].mult/added[3] ), .B(n11676), 
        .Y(n11675) );
  INVX1 U8593 ( .A(n11675), .Y(n11651) );
  INVX1 U8594 ( .A(\lamb/scale_ds1/genblk1[2].mult/added[1] ), .Y(n11652) );
  NAND2X1 U8595 ( .A(\lamb/scale_ds1/genblk1[2].mult/added[4] ), .B(
        \add_x_147/n1 ), .Y(n11552) );
  NAND3X1 U8596 ( .A(n11651), .B(n11652), .C(n11552), .Y(n11690) );
  INVX1 U8597 ( .A(\lamb/scale_ds1/genblk1[2].mult/added[2] ), .Y(n11674) );
  NAND3X1 U8598 ( .A(\lamb/scale_ds1/genblk1[2].mult/added[3] ), .B(
        \lamb/scale_ds1/genblk1[2].mult/added[4] ), .C(\add_x_147/n1 ), .Y(
        n11677) );
  AOI22X1 U8599 ( .A(n11553), .B(n11083), .C(n11674), .D(n10504), .Y(n11658)
         );
  AOI21X1 U8600 ( .A(\lamb/scale_ds1/genblk1[2].mult/added[4] ), .B(
        \add_x_147/n1 ), .C(\lamb/scale_ds1/genblk1[2].mult/added[3] ), .Y(
        n11650) );
  INVX1 U8601 ( .A(n10504), .Y(n11653) );
  NAND2X1 U8602 ( .A(\lamb/scale_ds1/genblk1[2].mult/added[2] ), .B(
        \lamb/scale_ds1/genblk1[2].mult/added[1] ), .Y(n11680) );
  OAI21X1 U8603 ( .A(n11653), .B(n11680), .C(n11554), .Y(n11654) );
  AOI21X1 U8604 ( .A(n11652), .B(n11166), .C(n11654), .Y(n11635) );
  AND2X1 U8605 ( .A(\lamb/scale_ts0/genblk1[1].mult/added[4] ), .B(
        \add_x_153/n1 ), .Y(n11555) );
  NAND2X1 U8606 ( .A(\lamb/scale_ts0/genblk1[1].mult/added[3] ), .B(n11555), 
        .Y(n11582) );
  INVX1 U8607 ( .A(n11582), .Y(n11556) );
  INVX1 U8608 ( .A(\lamb/scale_ts0/genblk1[1].mult/added[1] ), .Y(n11600) );
  NAND3X1 U8609 ( .A(n11556), .B(\lamb/scale_ts0/genblk1[1].mult/added[2] ), 
        .C(n11600), .Y(n11585) );
  NOR3X1 U8610 ( .A(\lamb/scale_ts0/genblk1[1].mult/added[3] ), .B(
        \lamb/scale_ts0/genblk1[1].mult/added[4] ), .C(\add_x_153/n1 ), .Y(
        n11581) );
  INVX1 U8611 ( .A(\lamb/scale_ts0/genblk1[1].mult/added[2] ), .Y(n11560) );
  AOI22X1 U8612 ( .A(\lamb/scale_ts0/genblk1[1].mult/added[2] ), .B(n11581), 
        .C(n11556), .D(n11560), .Y(n11617) );
  INVX1 U8613 ( .A(\lamb/scale_ts0/genblk1[1].mult/added[3] ), .Y(n11558) );
  NOR2X1 U8614 ( .A(\lamb/scale_ts0/genblk1[1].mult/added[4] ), .B(
        \add_x_153/n1 ), .Y(n11557) );
  AOI21X1 U8615 ( .A(\add_x_153/n1 ), .B(
        \lamb/scale_ts0/genblk1[1].mult/added[4] ), .C(n11557), .Y(n11559) );
  NAND2X1 U8616 ( .A(\lamb/scale_ts0/genblk1[1].mult/added[2] ), .B(n11619), 
        .Y(n11565) );
  NAND2X1 U8617 ( .A(\lamb/scale_ts0/genblk1[1].mult/added[3] ), .B(n10997), 
        .Y(n11580) );
  INVX1 U8618 ( .A(n11580), .Y(n11621) );
  NAND3X1 U8619 ( .A(n10443), .B(n11565), .C(n10965), .Y(n11567) );
  INVX1 U8620 ( .A(\lamb/scale_ts0/genblk1[1].mult/added[4] ), .Y(n11562) );
  AOI22X1 U8621 ( .A(\lamb/scale_ts0/genblk1[1].mult/added[4] ), .B(
        \lamb/scale_ts0/genblk1[1].mult/added[3] ), .C(\add_x_153/n1 ), .D(
        n11562), .Y(n11563) );
  OAI21X1 U8622 ( .A(\lamb/scale_ts0/genblk1[1].mult/added[3] ), .B(
        \add_x_153/n1 ), .C(n11563), .Y(n11583) );
  NAND2X1 U8623 ( .A(\lamb/scale_ts0/genblk1[1].mult/added[1] ), .B(n11581), 
        .Y(n11564) );
  AOI22X1 U8624 ( .A(\lamb/scale_ts0/genblk1[1].mult/added[1] ), .B(n11567), 
        .C(n10642), .D(n11566), .Y(n11569) );
  AOI21X1 U8625 ( .A(n13371), .B(n11127), .C(n13377), .Y(n13368) );
  NAND2X1 U8626 ( .A(n12293), .B(n13367), .Y(n13823) );
  AND2X1 U8627 ( .A(n11568), .B(n13823), .Y(n13378) );
  NAND2X1 U8628 ( .A(n13368), .B(n13378), .Y(n13385) );
  AOI21X1 U8629 ( .A(n11585), .B(n11569), .C(n10723), .Y(n11578) );
  MUX2X1 U8630 ( .B(n11571), .A(msg[51]), .S(n11570), .Y(n11572) );
  FAX1 U8631 ( .A(n11574), .B(n11573), .C(n11572), .YS(n11575) );
  FAX1 U8632 ( .A(n11577), .B(n11576), .C(n11575), .YS(n12671) );
  INVX1 U8633 ( .A(n12671), .Y(n12665) );
  HAX1 U8634 ( .A(n11578), .B(n12665), .YS(n13342) );
  INVX1 U8635 ( .A(n13342), .Y(n13347) );
  NAND2X1 U8636 ( .A(\lamb/scale_ts0/genblk1[1].mult/added[2] ), .B(n11600), 
        .Y(n11579) );
  OAI21X1 U8637 ( .A(n11580), .B(n11579), .C(n10443), .Y(n11602) );
  AOI21X1 U8638 ( .A(n11620), .B(n11582), .C(n11581), .Y(n11601) );
  NAND2X1 U8639 ( .A(n10954), .B(\lamb/scale_ts0/genblk1[1].mult/added[1] ), 
        .Y(n11584) );
  NAND3X1 U8640 ( .A(n11585), .B(n11077), .C(n11584), .Y(n11586) );
  OAI21X1 U8641 ( .A(n11602), .B(n11586), .C(n11622), .Y(n11599) );
  HAX1 U8642 ( .A(n11588), .B(n11587), .YS(n11589) );
  MUX2X1 U8643 ( .B(msg[1]), .A(n13815), .S(n11589), .Y(n12657) );
  INVX1 U8644 ( .A(n12657), .Y(n12658) );
  MUX2X1 U8645 ( .B(msg[2]), .A(n13811), .S(n11590), .Y(n11625) );
  HAX1 U8646 ( .A(n11105), .B(n11591), .YS(n11612) );
  MUX2X1 U8647 ( .B(n13711), .A(msg[29]), .S(n11593), .Y(n11594) );
  MUX2X1 U8648 ( .B(n11595), .A(msg[54]), .S(n11594), .Y(n11596) );
  FAX1 U8649 ( .A(n11625), .B(n11612), .C(n11596), .YS(n11597) );
  FAX1 U8650 ( .A(n11598), .B(n12658), .C(n11597), .YS(n12667) );
  AND2X1 U8651 ( .A(n13347), .B(n13349), .Y(n13341) );
  AOI22X1 U8652 ( .A(\lamb/scale_ts0/genblk1[1].mult/added[1] ), .B(n11077), 
        .C(n11619), .D(n11600), .Y(n11604) );
  INVX1 U8653 ( .A(n11602), .Y(n11603) );
  AOI21X1 U8654 ( .A(n11604), .B(n11603), .C(n10723), .Y(n11616) );
  HAX1 U8655 ( .A(n11145), .B(n11605), .YS(n11629) );
  INVX1 U8656 ( .A(n11606), .Y(n11609) );
  FAX1 U8657 ( .A(n11609), .B(n11608), .C(n11607), .YS(n11610) );
  FAX1 U8658 ( .A(msg[50]), .B(msg[53]), .C(n11610), .YS(n11611) );
  FAX1 U8659 ( .A(n11613), .B(n11612), .C(n11611), .YS(n11614) );
  FAX1 U8660 ( .A(n11615), .B(n11629), .C(n11614), .YS(n12659) );
  HAX1 U8661 ( .A(n11616), .B(n12659), .YS(n13350) );
  INVX1 U8662 ( .A(n13349), .Y(n12292) );
  INVX1 U8663 ( .A(n10443), .Y(n11618) );
  OAI21X1 U8664 ( .A(n11619), .B(n11618), .C(
        \lamb/scale_ts0/genblk1[1].mult/added[1] ), .Y(n11624) );
  AOI22X1 U8665 ( .A(\lamb/scale_ts0/genblk1[1].mult/added[2] ), .B(n10954), 
        .C(n11621), .D(n10642), .Y(n11623) );
  AOI21X1 U8666 ( .A(n11624), .B(n11623), .C(n10723), .Y(n11634) );
  MUX2X1 U8667 ( .B(n13729), .A(msg[22]), .S(n11625), .Y(n11630) );
  HAX1 U8668 ( .A(n11627), .B(n11156), .YS(n11628) );
  FAX1 U8669 ( .A(n11630), .B(n11629), .C(n11628), .YS(n11632) );
  FAX1 U8670 ( .A(n11633), .B(n11632), .C(n11631), .YS(n12670) );
  INVX1 U8671 ( .A(n12670), .Y(n12664) );
  HAX1 U8672 ( .A(n11634), .B(n12664), .YS(n13348) );
  AOI21X1 U8673 ( .A(n13350), .B(n10626), .C(n13348), .Y(n13340) );
  OAI21X1 U8674 ( .A(n11658), .B(n11635), .C(n11153), .Y(n11649) );
  OR2X1 U8675 ( .A(\add_x_143/n1 ), .B(
        \lamb/scale_ts1/genblk1[2].mult/added[4] ), .Y(n11641) );
  NAND2X1 U8676 ( .A(\lamb/scale_ts1/genblk1[2].mult/added[3] ), .B(n11641), 
        .Y(n11637) );
  INVX1 U8677 ( .A(\lamb/scale_ts1/genblk1[2].mult/added[3] ), .Y(n11640) );
  NAND2X1 U8678 ( .A(n11640), .B(n10397), .Y(n11636) );
  INVX1 U8679 ( .A(\lamb/scale_ts1/genblk1[2].mult/added[1] ), .Y(n11667) );
  NAND3X1 U8680 ( .A(\add_x_143/n1 ), .B(
        \lamb/scale_ts1/genblk1[2].mult/added[4] ), .C(
        \lamb/scale_ts1/genblk1[2].mult/added[3] ), .Y(n11644) );
  OAI21X1 U8681 ( .A(n11128), .B(n11667), .C(n11644), .Y(n11638) );
  OR2X1 U8682 ( .A(n11641), .B(\lamb/scale_ts1/genblk1[2].mult/added[3] ), .Y(
        n11643) );
  AND2X1 U8683 ( .A(\lamb/scale_ts1/genblk1[2].mult/added[2] ), .B(n11643), 
        .Y(n11668) );
  INVX1 U8684 ( .A(n11637), .Y(n11699) );
  AND2X1 U8685 ( .A(n11667), .B(n11699), .Y(n11661) );
  NAND2X1 U8686 ( .A(n11661), .B(n10397), .Y(n11702) );
  NAND2X1 U8687 ( .A(n11668), .B(n11702), .Y(n11659) );
  OAI21X1 U8688 ( .A(\lamb/scale_ts1/genblk1[2].mult/added[2] ), .B(n11638), 
        .C(n11659), .Y(n11663) );
  INVX1 U8689 ( .A(n11642), .Y(n11697) );
  INVX1 U8690 ( .A(n11643), .Y(n11645) );
  AND2X1 U8691 ( .A(\lamb/scale_ts1/genblk1[2].mult/added[2] ), .B(
        \lamb/scale_ts1/genblk1[2].mult/added[1] ), .Y(n11696) );
  OAI21X1 U8692 ( .A(n11645), .B(n11696), .C(n11644), .Y(n11662) );
  OAI21X1 U8693 ( .A(\lamb/scale_ts1/genblk1[2].mult/added[1] ), .B(n11697), 
        .C(n11662), .Y(n11647) );
  OAI21X1 U8694 ( .A(n13372), .B(n10851), .C(n11646), .Y(n13262) );
  INVX1 U8695 ( .A(n13262), .Y(n13273) );
  NOR2X1 U8696 ( .A(n12682), .B(n11709), .Y(n13256) );
  AOI21X1 U8697 ( .A(n13370), .B(n12682), .C(n13256), .Y(n13275) );
  INVX1 U8698 ( .A(n13275), .Y(n13269) );
  NAND2X1 U8699 ( .A(n13262), .B(n13269), .Y(n13260) );
  INVX1 U8700 ( .A(n13260), .Y(n13266) );
  AOI22X1 U8701 ( .A(n10851), .B(n12679), .C(n13377), .D(n12682), .Y(n13261)
         );
  OAI21X1 U8702 ( .A(n13266), .B(n13267), .C(n10471), .Y(n13263) );
  OAI21X1 U8703 ( .A(n11020), .B(n13263), .C(n12304), .Y(n11669) );
  AOI21X1 U8704 ( .A(n11663), .B(n11647), .C(n11669), .Y(n11648) );
  HAX1 U8705 ( .A(n11649), .B(n11648), .YS(n13877) );
  INVX1 U8706 ( .A(n13877), .Y(n13880) );
  AOI22X1 U8707 ( .A(\lamb/scale_ds1/genblk1[2].mult/added[1] ), .B(n10603), 
        .C(n11653), .D(n11652), .Y(n11656) );
  INVX1 U8708 ( .A(n11654), .Y(n11655) );
  NAND2X1 U8709 ( .A(n11656), .B(n11655), .Y(n11657) );
  OAI21X1 U8710 ( .A(n11658), .B(n11657), .C(n11153), .Y(n11666) );
  INVX1 U8711 ( .A(n11669), .Y(n11704) );
  INVX1 U8712 ( .A(n11659), .Y(n11660) );
  NAND3X1 U8713 ( .A(n11663), .B(n11662), .C(n11080), .Y(n11664) );
  NAND2X1 U8714 ( .A(n11704), .B(n11664), .Y(n11665) );
  HAX1 U8715 ( .A(n11666), .B(n11665), .YS(n13876) );
  AOI22X1 U8716 ( .A(\lamb/scale_ts1/genblk1[2].mult/added[1] ), .B(n11668), 
        .C(n11128), .D(n11667), .Y(n11698) );
  MUX2X1 U8717 ( .B(n11698), .A(\lamb/scale_ts1/genblk1[2].mult/added[2] ), 
        .S(n11697), .Y(n11671) );
  AOI21X1 U8718 ( .A(n11671), .B(n11080), .C(n11669), .Y(n11686) );
  AOI21X1 U8719 ( .A(n11675), .B(n11674), .C(n10911), .Y(n11687) );
  INVX1 U8720 ( .A(n11676), .Y(n11679) );
  NAND2X1 U8721 ( .A(n11166), .B(n10504), .Y(n11678) );
  AOI22X1 U8722 ( .A(n11679), .B(\lamb/scale_ds1/genblk1[2].mult/added[1] ), 
        .C(\lamb/scale_ds1/genblk1[2].mult/added[2] ), .D(n11678), .Y(n11683)
         );
  INVX1 U8723 ( .A(n10603), .Y(n11682) );
  INVX1 U8724 ( .A(n11680), .Y(n11681) );
  AOI22X1 U8725 ( .A(n11683), .B(n11682), .C(n11681), .D(n11166), .Y(n11684)
         );
  OAI21X1 U8726 ( .A(n11687), .B(n11684), .C(n11153), .Y(n11685) );
  HAX1 U8727 ( .A(n11686), .B(n11685), .YS(n13194) );
  INVX1 U8728 ( .A(n11687), .Y(n11692) );
  AOI22X1 U8729 ( .A(\lamb/scale_ds1/genblk1[2].mult/added[2] ), .B(n10603), 
        .C(\lamb/scale_ds1/genblk1[2].mult/added[1] ), .D(n11688), .Y(n11691)
         );
  NAND3X1 U8730 ( .A(n11692), .B(n11691), .C(n11083), .Y(n11694) );
  NAND2X1 U8731 ( .A(n11694), .B(n11153), .Y(n11706) );
  AOI22X1 U8732 ( .A(\lamb/scale_ts1/genblk1[2].mult/added[1] ), .B(n11697), 
        .C(n11695), .D(n11696), .Y(n11701) );
  OAI21X1 U8733 ( .A(\lamb/scale_ts1/genblk1[2].mult/added[2] ), .B(n11699), 
        .C(n11698), .Y(n11700) );
  NAND3X1 U8734 ( .A(n11702), .B(n11701), .C(n11700), .Y(n11703) );
  HAX1 U8735 ( .A(n11706), .B(n10972), .YS(n13195) );
  INVX1 U8736 ( .A(n13195), .Y(n13879) );
  NOR3X1 U8737 ( .A(n13880), .B(n13876), .C(n11054), .Y(n11774) );
  AOI21X1 U8738 ( .A(n11707), .B(n11739), .C(n11774), .Y(n11729) );
  NAND2X1 U8739 ( .A(n13337), .B(n10809), .Y(n11708) );
  OAI21X1 U8740 ( .A(n11709), .B(n10635), .C(n11708), .Y(n13158) );
  INVX1 U8741 ( .A(n13830), .Y(n13333) );
  NAND2X1 U8742 ( .A(n13333), .B(n10809), .Y(n11710) );
  OAI21X1 U8743 ( .A(n11711), .B(n10635), .C(n11710), .Y(n13157) );
  INVX1 U8744 ( .A(n10440), .Y(n12699) );
  NAND3X1 U8745 ( .A(n13229), .B(n12699), .C(n11712), .Y(n12700) );
  OAI21X1 U8746 ( .A(n13235), .B(n13336), .C(n12700), .Y(n13154) );
  NAND2X1 U8747 ( .A(n13157), .B(n13154), .Y(n11715) );
  OAI21X1 U8748 ( .A(n13834), .B(n11713), .C(n11714), .Y(n12511) );
  INVX1 U8749 ( .A(n12511), .Y(n13161) );
  AOI21X1 U8750 ( .A(n13158), .B(n11715), .C(n13161), .Y(n13155) );
  INVX1 U8751 ( .A(n13154), .Y(n13167) );
  NAND2X1 U8752 ( .A(n13161), .B(n13167), .Y(n13168) );
  INVX1 U8753 ( .A(n13158), .Y(n13160) );
  INVX1 U8754 ( .A(n12215), .Y(n12438) );
  AOI21X1 U8755 ( .A(n11023), .B(n13169), .C(n12438), .Y(n11779) );
  OR2X1 U8756 ( .A(\add_x_129/n1 ), .B(
        \lamb/scale_ts2/genblk1[3].mult/added[4] ), .Y(n11717) );
  NAND2X1 U8757 ( .A(\lamb/scale_ts2/genblk1[3].mult/added[3] ), .B(n11717), 
        .Y(n11723) );
  INVX1 U8758 ( .A(n11723), .Y(n11716) );
  INVX1 U8759 ( .A(\lamb/scale_ts2/genblk1[3].mult/added[1] ), .Y(n11751) );
  NAND3X1 U8760 ( .A(n11716), .B(n11751), .C(n10510), .Y(n11747) );
  INVX1 U8761 ( .A(\lamb/scale_ts2/genblk1[3].mult/added[3] ), .Y(n11722) );
  INVX1 U8762 ( .A(n11750), .Y(n11720) );
  INVX1 U8763 ( .A(\add_x_129/n1 ), .Y(n11718) );
  AOI22X1 U8764 ( .A(\add_x_129/n1 ), .B(
        \lamb/scale_ts2/genblk1[3].mult/added[4] ), .C(
        \lamb/scale_ts2/genblk1[3].mult/added[3] ), .D(n11718), .Y(n11719) );
  AOI21X1 U8765 ( .A(\lamb/scale_ts2/genblk1[3].mult/added[4] ), .B(
        \lamb/scale_ts2/genblk1[3].mult/added[3] ), .C(n11719), .Y(n11754) );
  AOI22X1 U8766 ( .A(\lamb/scale_ts2/genblk1[3].mult/added[1] ), .B(n11720), 
        .C(\lamb/scale_ts2/genblk1[3].mult/added[2] ), .D(n10637), .Y(n11726)
         );
  NAND2X1 U8767 ( .A(n11722), .B(n10510), .Y(n11724) );
  INVX1 U8768 ( .A(\lamb/scale_ts2/genblk1[3].mult/added[2] ), .Y(n11743) );
  MUX2X1 U8769 ( .B(n11724), .A(n11723), .S(n11743), .Y(n11725) );
  NAND3X1 U8770 ( .A(n11747), .B(n11726), .C(n11002), .Y(n11727) );
  NAND2X1 U8771 ( .A(n10679), .B(n11727), .Y(n11728) );
  HAX1 U8772 ( .A(n11729), .B(n11728), .YS(n13101) );
  INVX1 U8773 ( .A(n13101), .Y(n13099) );
  NAND3X1 U8774 ( .A(\add_x_129/n1 ), .B(
        \lamb/scale_ts2/genblk1[3].mult/added[4] ), .C(
        \lamb/scale_ts2/genblk1[3].mult/added[3] ), .Y(n11745) );
  NAND2X1 U8775 ( .A(n11750), .B(n10386), .Y(n11731) );
  NOR3X1 U8776 ( .A(\add_x_129/n1 ), .B(
        \lamb/scale_ts2/genblk1[3].mult/added[4] ), .C(
        \lamb/scale_ts2/genblk1[3].mult/added[3] ), .Y(n11746) );
  AOI22X1 U8777 ( .A(\lamb/scale_ts2/genblk1[3].mult/added[2] ), .B(n11731), 
        .C(\lamb/scale_ts2/genblk1[3].mult/added[1] ), .D(n11746), .Y(n11733)
         );
  INVX1 U8778 ( .A(n10637), .Y(n11732) );
  AOI22X1 U8779 ( .A(\lamb/scale_ts2/genblk1[3].mult/added[1] ), .B(
        \lamb/scale_ts2/genblk1[3].mult/added[2] ), .C(n11733), .D(n11732), 
        .Y(n11752) );
  OAI21X1 U8780 ( .A(n11730), .B(n10422), .C(n10679), .Y(n11742) );
  INVX1 U8781 ( .A(n11734), .Y(n11735) );
  NAND3X1 U8782 ( .A(n11759), .B(n11736), .C(n11735), .Y(n11765) );
  NAND2X1 U8783 ( .A(n11761), .B(\lamb/scale_ds2/genblk1[3].mult/added[1] ), 
        .Y(n11737) );
  AOI22X1 U8784 ( .A(\lamb/scale_ds2/genblk1[3].mult/added[2] ), .B(n11773), 
        .C(n10427), .D(n11738), .Y(n11740) );
  AOI21X1 U8785 ( .A(n11740), .B(n11739), .C(n11774), .Y(n11741) );
  XNOR2X1 U8786 ( .A(n11742), .B(n10387), .Y(n13100) );
  OAI21X1 U8787 ( .A(n10926), .B(n11746), .C(n10386), .Y(n11778) );
  INVX1 U8788 ( .A(n10386), .Y(n11753) );
  INVX1 U8789 ( .A(n11746), .Y(n11748) );
  NAND3X1 U8790 ( .A(n11748), .B(n11747), .C(
        \lamb/scale_ts2/genblk1[3].mult/added[2] ), .Y(n11749) );
  OAI21X1 U8791 ( .A(\lamb/scale_ts2/genblk1[3].mult/added[2] ), .B(n11753), 
        .C(n11749), .Y(n11782) );
  NAND2X1 U8792 ( .A(n11751), .B(n11750), .Y(n11777) );
  AOI22X1 U8793 ( .A(n10637), .B(n11777), .C(n11753), .D(n10422), .Y(n11755)
         );
  NAND3X1 U8794 ( .A(n11778), .B(n11782), .C(n11755), .Y(n11756) );
  NAND2X1 U8795 ( .A(n10679), .B(n11756), .Y(n11770) );
  AOI22X1 U8796 ( .A(\lamb/scale_ds2/genblk1[3].mult/added[3] ), .B(n11759), 
        .C(n11168), .D(n10427), .Y(n11771) );
  AOI21X1 U8797 ( .A(n10947), .B(\lamb/scale_ds2/genblk1[3].mult/added[1] ), 
        .C(n11771), .Y(n11766) );
  NOR2X1 U8798 ( .A(n11760), .B(n11151), .Y(n11764) );
  NAND3X1 U8799 ( .A(\lamb/scale_ds2/genblk1[3].mult/added[2] ), .B(n11762), 
        .C(n11168), .Y(n11763) );
  OAI21X1 U8800 ( .A(\lamb/scale_ds2/genblk1[3].mult/added[2] ), .B(n11764), 
        .C(n11763), .Y(n11776) );
  NAND3X1 U8801 ( .A(n11766), .B(n11765), .C(n11776), .Y(n11768) );
  INVX1 U8802 ( .A(n11774), .Y(n11767) );
  HAX1 U8803 ( .A(n11770), .B(n10970), .YS(n13097) );
  INVX1 U8804 ( .A(n13097), .Y(n13091) );
  INVX1 U8805 ( .A(n11771), .Y(n11772) );
  OAI21X1 U8806 ( .A(\lamb/scale_ds2/genblk1[3].mult/added[1] ), .B(n11773), 
        .C(n11772), .Y(n11775) );
  AOI21X1 U8807 ( .A(n11776), .B(n11775), .C(n11774), .Y(n11784) );
  NAND2X1 U8808 ( .A(n11778), .B(n11777), .Y(n11781) );
  INVX1 U8809 ( .A(n10679), .Y(n11780) );
  AOI21X1 U8810 ( .A(n11782), .B(n11781), .C(n11780), .Y(n11783) );
  HAX1 U8811 ( .A(n11784), .B(n10969), .YS(n13092) );
  INVX1 U8812 ( .A(n13092), .Y(n13098) );
  NAND3X1 U8813 ( .A(n11076), .B(n13091), .C(n13098), .Y(n12514) );
  OAI21X1 U8814 ( .A(n10809), .B(n13841), .C(n10676), .Y(n11785) );
  AOI21X1 U8815 ( .A(n10799), .B(n13841), .C(n11785), .Y(n11989) );
  INVX1 U8816 ( .A(\lamb/scale_bs3/genblk1[0].mult/added[3] ), .Y(n11788) );
  INVX1 U8817 ( .A(\lamb/scale_bs3/genblk1[0].mult/added[1] ), .Y(n11786) );
  NAND3X1 U8818 ( .A(\lamb/scale_bs3/genblk1[0].mult/added[2] ), .B(n11122), 
        .C(n11786), .Y(n11931) );
  NAND2X1 U8819 ( .A(\lamb/scale_bs3/genblk1[0].mult/added[2] ), .B(
        \lamb/scale_bs3/genblk1[0].mult/added[1] ), .Y(n11929) );
  INVX1 U8820 ( .A(n11929), .Y(n11983) );
  NOR3X1 U8821 ( .A(\lamb/scale_bs3/genblk1[0].mult/added[4] ), .B(
        \add_x_125/n1 ), .C(\lamb/scale_bs3/genblk1[0].mult/added[3] ), .Y(
        n11808) );
  AOI21X1 U8822 ( .A(n11983), .B(n11789), .C(n11808), .Y(n11807) );
  NOR2X1 U8823 ( .A(\lamb/scale_bs3/genblk1[0].mult/added[4] ), .B(
        \add_x_125/n1 ), .Y(n11920) );
  INVX1 U8824 ( .A(n11920), .Y(n11806) );
  NAND3X1 U8825 ( .A(n11927), .B(n11786), .C(n10641), .Y(n11987) );
  NAND2X1 U8826 ( .A(n11788), .B(n10641), .Y(n11805) );
  NAND2X1 U8827 ( .A(n11805), .B(n11114), .Y(n11921) );
  INVX1 U8828 ( .A(n11921), .Y(n11982) );
  AOI21X1 U8829 ( .A(n11982), .B(\lamb/scale_bs3/genblk1[0].mult/added[1] ), 
        .C(n11122), .Y(n11790) );
  INVX1 U8830 ( .A(\lamb/scale_bs3/genblk1[0].mult/added[2] ), .Y(n11923) );
  AOI22X1 U8831 ( .A(\lamb/scale_bs3/genblk1[0].mult/added[2] ), .B(n11987), 
        .C(n11790), .D(n11923), .Y(n11811) );
  INVX1 U8832 ( .A(n11811), .Y(n11791) );
  NAND3X1 U8833 ( .A(n11931), .B(n10421), .C(n11791), .Y(n11792) );
  NAND2X1 U8834 ( .A(n10675), .B(n11792), .Y(n11793) );
  HAX1 U8835 ( .A(n11794), .B(n11793), .YS(n12161) );
  INVX1 U8836 ( .A(n12161), .Y(n12035) );
  OR2X1 U8837 ( .A(\lamb/scale_ls3/genblk1[2].mult/added[4] ), .B(
        \add_x_126/n1 ), .Y(n11944) );
  AOI21X1 U8838 ( .A(\lamb/scale_ls3/genblk1[2].mult/added[2] ), .B(
        \lamb/scale_ls3/genblk1[2].mult/added[1] ), .C(n10441), .Y(n11940) );
  INVX1 U8839 ( .A(\lamb/scale_ls3/genblk1[2].mult/added[2] ), .Y(n11943) );
  INVX1 U8840 ( .A(\lamb/scale_ls3/genblk1[2].mult/added[3] ), .Y(n11891) );
  NAND2X1 U8841 ( .A(n11891), .B(n11194), .Y(n11795) );
  NAND2X1 U8842 ( .A(n11795), .B(n10441), .Y(n11892) );
  NAND3X1 U8843 ( .A(n11944), .B(n11891), .C(n11194), .Y(n11890) );
  OR2X1 U8844 ( .A(\lamb/scale_ls3/genblk1[2].mult/added[3] ), .B(n11944), .Y(
        n11894) );
  INVX1 U8845 ( .A(n11894), .Y(n11797) );
  NAND2X1 U8846 ( .A(\lamb/scale_ls3/genblk1[2].mult/added[3] ), .B(n11937), 
        .Y(n11945) );
  INVX1 U8847 ( .A(n11945), .Y(n11796) );
  AOI22X1 U8848 ( .A(\lamb/scale_ls3/genblk1[2].mult/added[2] ), .B(n11797), 
        .C(n11796), .D(n11943), .Y(n11951) );
  INVX1 U8849 ( .A(\lamb/scale_ls3/genblk1[2].mult/added[1] ), .Y(n11941) );
  AOI21X1 U8850 ( .A(n11890), .B(n11951), .C(n11941), .Y(n11798) );
  INVX1 U8851 ( .A(n11798), .Y(n11799) );
  OAI21X1 U8852 ( .A(n11943), .B(n11892), .C(n11799), .Y(n11800) );
  AOI21X1 U8853 ( .A(n11940), .B(n11194), .C(n11800), .Y(n12058) );
  XNOR2X1 U8854 ( .A(n12035), .B(n10840), .Y(n12084) );
  NOR3X1 U8855 ( .A(\lamb/scale_ls3/genblk1[0].mult/added[3] ), .B(n11542), 
        .C(n11910), .Y(n11991) );
  AOI22X1 U8856 ( .A(\lamb/scale_ls3/genblk1[0].mult/added[1] ), .B(n11051), 
        .C(n11991), .D(n11801), .Y(n11803) );
  AOI21X1 U8857 ( .A(n11804), .B(n11803), .C(n11995), .Y(n11813) );
  INVX1 U8858 ( .A(n11805), .Y(n11925) );
  NAND2X1 U8859 ( .A(n11925), .B(n11806), .Y(n11919) );
  AOI22X1 U8860 ( .A(\lamb/scale_bs3/genblk1[0].mult/added[2] ), .B(n11808), 
        .C(\lamb/scale_bs3/genblk1[0].mult/added[1] ), .D(n10421), .Y(n11809)
         );
  OAI21X1 U8861 ( .A(n11983), .B(n11919), .C(n11809), .Y(n11810) );
  OAI21X1 U8862 ( .A(n11811), .B(n11810), .C(n10675), .Y(n11812) );
  HAX1 U8863 ( .A(n11813), .B(n11812), .YS(n12090) );
  NAND3X1 U8864 ( .A(\lamb/scale_ls3/genblk1[1].mult/added[3] ), .B(
        \add_x_127/n1 ), .C(\lamb/scale_ls3/genblk1[1].mult/added[4] ), .Y(
        n11815) );
  INVX1 U8865 ( .A(n11815), .Y(n11820) );
  INVX1 U8866 ( .A(\lamb/scale_ls3/genblk1[1].mult/added[1] ), .Y(n11817) );
  NAND3X1 U8867 ( .A(n11820), .B(\lamb/scale_ls3/genblk1[1].mult/added[2] ), 
        .C(n11817), .Y(n11966) );
  OR2X1 U8868 ( .A(\add_x_127/n1 ), .B(
        \lamb/scale_ls3/genblk1[1].mult/added[4] ), .Y(n11877) );
  AOI21X1 U8869 ( .A(\add_x_127/n1 ), .B(
        \lamb/scale_ls3/genblk1[1].mult/added[4] ), .C(
        \lamb/scale_ls3/genblk1[1].mult/added[3] ), .Y(n11899) );
  AOI21X1 U8870 ( .A(\lamb/scale_ls3/genblk1[1].mult/added[3] ), .B(n11877), 
        .C(n10654), .Y(n11876) );
  INVX1 U8871 ( .A(n11876), .Y(n11961) );
  NAND2X1 U8872 ( .A(\lamb/scale_ls3/genblk1[1].mult/added[3] ), .B(n11877), 
        .Y(n11814) );
  AOI21X1 U8873 ( .A(\add_x_127/n1 ), .B(
        \lamb/scale_ls3/genblk1[1].mult/added[4] ), .C(n11814), .Y(n11955) );
  INVX1 U8874 ( .A(\lamb/scale_ls3/genblk1[1].mult/added[2] ), .Y(n11954) );
  NOR2X1 U8875 ( .A(n11954), .B(\lamb/scale_ls3/genblk1[1].mult/added[1] ), 
        .Y(n11816) );
  NOR2X1 U8876 ( .A(n11877), .B(\lamb/scale_ls3/genblk1[1].mult/added[3] ), 
        .Y(n11958) );
  INVX1 U8877 ( .A(n11958), .Y(n11819) );
  AOI22X1 U8878 ( .A(\lamb/scale_ls3/genblk1[1].mult/added[2] ), .B(n11819), 
        .C(n11815), .D(n11954), .Y(n11953) );
  OAI21X1 U8879 ( .A(n11817), .B(n11961), .C(n11004), .Y(n11818) );
  INVX1 U8880 ( .A(n11818), .Y(n11822) );
  OAI21X1 U8881 ( .A(n11143), .B(n11820), .C(n11819), .Y(n11821) );
  INVX1 U8882 ( .A(n11821), .Y(n11898) );
  NAND3X1 U8883 ( .A(n11966), .B(n11822), .C(n11898), .Y(n11862) );
  AOI21X1 U8884 ( .A(\add_x_140/n1 ), .B(
        \lamb/scale_ls2/genblk1[1].mult/added[4] ), .C(
        \lamb/scale_ls2/genblk1[1].mult/added[3] ), .Y(n11846) );
  OR2X1 U8885 ( .A(\add_x_140/n1 ), .B(
        \lamb/scale_ls2/genblk1[1].mult/added[4] ), .Y(n11823) );
  AND2X1 U8886 ( .A(n10555), .B(n11823), .Y(n11856) );
  INVX1 U8887 ( .A(n10555), .Y(n11838) );
  NAND2X1 U8888 ( .A(n10752), .B(n11838), .Y(n11853) );
  INVX1 U8889 ( .A(\lamb/scale_ls2/genblk1[1].mult/added[2] ), .Y(n11832) );
  AND2X1 U8890 ( .A(\add_x_140/n1 ), .B(
        \lamb/scale_ls2/genblk1[1].mult/added[4] ), .Y(n11830) );
  OR2X1 U8891 ( .A(n11832), .B(n10643), .Y(n11841) );
  NOR3X1 U8892 ( .A(\lamb/scale_ls2/genblk1[1].mult/added[3] ), .B(
        \add_x_140/n1 ), .C(\lamb/scale_ls2/genblk1[1].mult/added[4] ), .Y(
        n11836) );
  NAND2X1 U8893 ( .A(n11836), .B(\lamb/scale_ls2/genblk1[1].mult/added[1] ), 
        .Y(n11824) );
  NAND3X1 U8894 ( .A(n11853), .B(n11841), .C(n11824), .Y(n11825) );
  AOI22X1 U8895 ( .A(\lamb/scale_ls2/genblk1[1].mult/added[2] ), .B(n11856), 
        .C(n11001), .D(n11825), .Y(n11827) );
  NOR2X1 U8896 ( .A(n11832), .B(n11836), .Y(n11833) );
  INVX1 U8897 ( .A(n11833), .Y(n11826) );
  NAND3X1 U8898 ( .A(\lamb/scale_ls2/genblk1[1].mult/added[1] ), .B(n11826), 
        .C(n11086), .Y(n11858) );
  AOI21X1 U8899 ( .A(n11827), .B(n11858), .C(n10799), .Y(n11829) );
  INVX1 U8900 ( .A(n13855), .Y(n13858) );
  NAND2X1 U8901 ( .A(n10809), .B(n13858), .Y(n11828) );
  HAX1 U8902 ( .A(n11829), .B(n11828), .YS(n13123) );
  INVX1 U8903 ( .A(n13123), .Y(n13119) );
  NOR3X1 U8904 ( .A(n10752), .B(\lamb/scale_ls2/genblk1[1].mult/added[1] ), 
        .C(n11830), .Y(n11831) );
  INVX1 U8905 ( .A(n11831), .Y(n11852) );
  AOI22X1 U8906 ( .A(n11833), .B(n11852), .C(n11832), .D(n10643), .Y(n11849)
         );
  OAI21X1 U8907 ( .A(n11834), .B(n11836), .C(n10643), .Y(n11845) );
  NAND3X1 U8908 ( .A(n11838), .B(\lamb/scale_ls2/genblk1[1].mult/added[1] ), 
        .C(n10752), .Y(n11839) );
  AND2X1 U8909 ( .A(n11845), .B(n11839), .Y(n11840) );
  OAI21X1 U8910 ( .A(\lamb/scale_ls2/genblk1[1].mult/added[1] ), .B(n11841), 
        .C(n11840), .Y(n11842) );
  OAI21X1 U8911 ( .A(n11849), .B(n11842), .C(n11857), .Y(n11844) );
  NAND2X1 U8912 ( .A(n10809), .B(n13846), .Y(n11843) );
  HAX1 U8913 ( .A(n11844), .B(n11843), .YS(n13122) );
  OR2X1 U8914 ( .A(n13119), .B(n13122), .Y(n13864) );
  NAND2X1 U8915 ( .A(n13119), .B(n13122), .Y(n13115) );
  INVX1 U8916 ( .A(n13115), .Y(n13117) );
  OAI21X1 U8917 ( .A(\lamb/scale_ls2/genblk1[1].mult/added[1] ), .B(n10555), 
        .C(n11845), .Y(n11847) );
  INVX1 U8918 ( .A(n11847), .Y(n11848) );
  OAI21X1 U8919 ( .A(n11849), .B(n11848), .C(n11857), .Y(n11851) );
  XNOR2X1 U8920 ( .A(n11851), .B(n10389), .Y(n13121) );
  NAND2X1 U8921 ( .A(n11853), .B(n11852), .Y(n11854) );
  AOI22X1 U8922 ( .A(\lamb/scale_ls2/genblk1[1].mult/added[1] ), .B(n11856), 
        .C(n11086), .D(n11854), .Y(n11859) );
  AOI21X1 U8923 ( .A(n11859), .B(n11858), .C(n10799), .Y(n11861) );
  NAND2X1 U8924 ( .A(n10809), .B(n13857), .Y(n11860) );
  HAX1 U8925 ( .A(n11861), .B(n11860), .YS(n13116) );
  OAI21X1 U8926 ( .A(n13117), .B(n13121), .C(n13116), .Y(n13863) );
  OR2X1 U8927 ( .A(n13864), .B(n13863), .Y(n11878) );
  INVX1 U8928 ( .A(n10462), .Y(n11974) );
  INVX1 U8929 ( .A(\lamb/scale_bs3/genblk1[1].mult/added[3] ), .Y(n11865) );
  INVX1 U8930 ( .A(\lamb/scale_bs3/genblk1[1].mult/added[1] ), .Y(n11866) );
  AOI22X1 U8931 ( .A(\lamb/scale_bs3/genblk1[1].mult/added[1] ), .B(
        \lamb/scale_bs3/genblk1[1].mult/added[2] ), .C(n11865), .D(n11866), 
        .Y(n11864) );
  NAND2X1 U8932 ( .A(\add_x_124/n1 ), .B(
        \lamb/scale_bs3/genblk1[1].mult/added[4] ), .Y(n11863) );
  NAND2X1 U8933 ( .A(n10731), .B(n11865), .Y(n11868) );
  NAND3X1 U8934 ( .A(\lamb/scale_bs3/genblk1[1].mult/added[2] ), .B(n11885), 
        .C(n11868), .Y(n11973) );
  NAND3X1 U8935 ( .A(\add_x_124/n1 ), .B(
        \lamb/scale_bs3/genblk1[1].mult/added[4] ), .C(
        \lamb/scale_bs3/genblk1[1].mult/added[3] ), .Y(n11869) );
  INVX1 U8936 ( .A(n11869), .Y(n11867) );
  OR2X1 U8937 ( .A(\lamb/scale_bs3/genblk1[1].mult/added[2] ), .B(n11867), .Y(
        n11881) );
  NAND2X1 U8938 ( .A(n11973), .B(n11881), .Y(n11906) );
  AOI21X1 U8939 ( .A(\lamb/scale_bs3/genblk1[1].mult/added[4] ), .B(
        \add_x_124/n1 ), .C(\lamb/scale_bs3/genblk1[1].mult/added[3] ), .Y(
        n11903) );
  INVX1 U8940 ( .A(n11903), .Y(n11883) );
  OAI21X1 U8941 ( .A(n11865), .B(n10731), .C(n11883), .Y(n11970) );
  INVX1 U8942 ( .A(n11970), .Y(n11884) );
  AOI22X1 U8943 ( .A(\lamb/scale_bs3/genblk1[1].mult/added[1] ), .B(n11884), 
        .C(n11867), .D(n11866), .Y(n11872) );
  AND2X1 U8944 ( .A(\lamb/scale_bs3/genblk1[1].mult/added[2] ), .B(
        \lamb/scale_bs3/genblk1[1].mult/added[1] ), .Y(n11871) );
  INVX1 U8945 ( .A(n11868), .Y(n11870) );
  OAI21X1 U8946 ( .A(n11871), .B(n11870), .C(n11869), .Y(n11902) );
  NAND3X1 U8947 ( .A(n11906), .B(n10933), .C(n11902), .Y(n11873) );
  NAND2X1 U8948 ( .A(n11974), .B(n11873), .Y(n11874) );
  HAX1 U8949 ( .A(n10979), .B(n11874), .YS(n13429) );
  INVX1 U8950 ( .A(n13429), .Y(n13478) );
  HAX1 U8951 ( .A(n12090), .B(n13478), .YS(n12144) );
  AOI22X1 U8952 ( .A(\lamb/scale_ls3/genblk1[1].mult/added[2] ), .B(n11876), 
        .C(n10507), .D(n11143), .Y(n11880) );
  AND2X1 U8953 ( .A(n10654), .B(n11877), .Y(n11952) );
  OAI21X1 U8954 ( .A(n11952), .B(n11953), .C(
        \lamb/scale_ls3/genblk1[1].mult/added[1] ), .Y(n11879) );
  INVX1 U8955 ( .A(n11878), .Y(n11965) );
  AOI21X1 U8956 ( .A(n11880), .B(n11879), .C(n11965), .Y(n11888) );
  NAND2X1 U8957 ( .A(n11881), .B(\lamb/scale_bs3/genblk1[1].mult/added[1] ), 
        .Y(n11882) );
  AOI21X1 U8958 ( .A(\lamb/scale_bs3/genblk1[1].mult/added[2] ), .B(n11883), 
        .C(n11882), .Y(n11971) );
  AOI21X1 U8959 ( .A(\lamb/scale_bs3/genblk1[1].mult/added[2] ), .B(n11884), 
        .C(n11971), .Y(n11886) );
  AOI21X1 U8960 ( .A(n11886), .B(n11885), .C(n10462), .Y(n11887) );
  HAX1 U8961 ( .A(n11888), .B(n11887), .YS(n13436) );
  NAND2X1 U8962 ( .A(n11937), .B(n11941), .Y(n11889) );
  NAND2X1 U8963 ( .A(n11890), .B(n11889), .Y(n11897) );
  OAI21X1 U8964 ( .A(n11891), .B(\lamb/scale_ls3/genblk1[2].mult/added[2] ), 
        .C(n11944), .Y(n11942) );
  INVX1 U8965 ( .A(n11942), .Y(n11893) );
  OAI21X1 U8966 ( .A(n11893), .B(n11941), .C(n11892), .Y(n11896) );
  NAND3X1 U8967 ( .A(\lamb/scale_ls3/genblk1[2].mult/added[2] ), .B(
        \lamb/scale_ls3/genblk1[2].mult/added[1] ), .C(n11894), .Y(n11895) );
  AOI22X1 U8968 ( .A(\lamb/scale_ls3/genblk1[2].mult/added[2] ), .B(n11897), 
        .C(n11896), .D(n11895), .Y(n12071) );
  HAX1 U8969 ( .A(n10842), .B(n12161), .YS(n12101) );
  OAI21X1 U8970 ( .A(\lamb/scale_ls3/genblk1[1].mult/added[1] ), .B(n10654), 
        .C(n11898), .Y(n11900) );
  AOI21X1 U8971 ( .A(n11004), .B(n11900), .C(n11965), .Y(n11908) );
  OAI21X1 U8972 ( .A(\lamb/scale_bs3/genblk1[1].mult/added[1] ), .B(n11903), 
        .C(n11902), .Y(n11905) );
  AOI21X1 U8973 ( .A(n11906), .B(n11905), .C(n10462), .Y(n11907) );
  HAX1 U8974 ( .A(n11908), .B(n11907), .YS(n13458) );
  NAND2X1 U8975 ( .A(n13458), .B(n13478), .Y(n13431) );
  NOR2X1 U8976 ( .A(n13478), .B(n13458), .Y(n13438) );
  INVX1 U8977 ( .A(n13438), .Y(n11909) );
  XNOR2X1 U8978 ( .A(n12035), .B(n12090), .Y(n12045) );
  XNOR2X1 U8979 ( .A(n11196), .B(n12045), .Y(n12080) );
  AOI21X1 U8980 ( .A(n11910), .B(\lamb/scale_ls3/genblk1[0].mult/added[1] ), 
        .C(n10588), .Y(n11913) );
  AOI21X1 U8981 ( .A(\lamb/scale_ls3/genblk1[0].mult/added[3] ), .B(
        \lamb/scale_ls3/genblk1[0].mult/added[2] ), .C(n11911), .Y(n11912) );
  OAI21X1 U8982 ( .A(\lamb/scale_ls3/genblk1[0].mult/added[3] ), .B(
        \lamb/scale_ls3/genblk1[0].mult/added[2] ), .C(n11912), .Y(n11994) );
  OAI21X1 U8983 ( .A(\lamb/scale_ls3/genblk1[0].mult/added[2] ), .B(n11913), 
        .C(n11994), .Y(n11918) );
  OAI21X1 U8984 ( .A(n11914), .B(n11991), .C(
        \lamb/scale_ls3/genblk1[0].mult/added[2] ), .Y(n11916) );
  AOI21X1 U8985 ( .A(n11916), .B(n11915), .C(
        \lamb/scale_ls3/genblk1[0].mult/added[1] ), .Y(n11917) );
  OAI21X1 U8986 ( .A(n11918), .B(n11917), .C(n10677), .Y(n11934) );
  INVX1 U8987 ( .A(n11919), .Y(n11981) );
  AOI22X1 U8988 ( .A(\lamb/scale_bs3/genblk1[0].mult/added[2] ), .B(n11981), 
        .C(\lamb/scale_bs3/genblk1[0].mult/added[1] ), .D(n11920), .Y(n11922)
         );
  NAND2X1 U8989 ( .A(n11922), .B(n11921), .Y(n11928) );
  NAND2X1 U8990 ( .A(\lamb/scale_bs3/genblk1[0].mult/added[1] ), .B(n11923), 
        .Y(n11979) );
  AOI22X1 U8991 ( .A(n11983), .B(n11925), .C(n11982), .D(n10942), .Y(n11926)
         );
  OAI21X1 U8992 ( .A(n11114), .B(n11979), .C(n11926), .Y(n11984) );
  AOI21X1 U8993 ( .A(n11929), .B(n11928), .C(n11984), .Y(n11932) );
  INVX1 U8994 ( .A(n10675), .Y(n11930) );
  AOI21X1 U8995 ( .A(n11932), .B(n11931), .C(n11930), .Y(n11933) );
  XNOR2X1 U8996 ( .A(n11934), .B(n10388), .Y(n12109) );
  AND2X1 U8997 ( .A(n11944), .B(n11943), .Y(n11938) );
  INVX1 U8998 ( .A(n10441), .Y(n11936) );
  AOI21X1 U8999 ( .A(n11938), .B(n11194), .C(n11936), .Y(n11939) );
  AOI22X1 U9000 ( .A(\lamb/scale_ls3/genblk1[2].mult/added[2] ), .B(n11940), 
        .C(\lamb/scale_ls3/genblk1[2].mult/added[1] ), .D(n11939), .Y(n11950)
         );
  OAI21X1 U9001 ( .A(n11937), .B(n11942), .C(n11941), .Y(n11948) );
  OAI21X1 U9002 ( .A(\lamb/scale_ls3/genblk1[2].mult/added[3] ), .B(n11944), 
        .C(n11943), .Y(n11946) );
  NAND3X1 U9003 ( .A(\lamb/scale_ls3/genblk1[2].mult/added[1] ), .B(n11946), 
        .C(n11945), .Y(n11947) );
  AOI21X1 U9004 ( .A(n11948), .B(n11947), .C(n11223), .Y(n12073) );
  NAND3X1 U9005 ( .A(n10840), .B(n10842), .C(n10843), .Y(n11949) );
  HAX1 U9006 ( .A(n12109), .B(n12132), .YS(n12037) );
  INVX1 U9007 ( .A(n12037), .Y(n12164) );
  NAND2X1 U9008 ( .A(\lamb/scale_ls3/genblk1[1].mult/added[2] ), .B(n11952), 
        .Y(n11960) );
  INVX1 U9009 ( .A(n11953), .Y(n11957) );
  NAND2X1 U9010 ( .A(n10507), .B(n11954), .Y(n11956) );
  NAND3X1 U9011 ( .A(n11960), .B(n11957), .C(n11956), .Y(n11964) );
  NAND2X1 U9012 ( .A(\lamb/scale_ls3/genblk1[1].mult/added[1] ), .B(n11958), 
        .Y(n11959) );
  NAND3X1 U9013 ( .A(n11961), .B(n11960), .C(n11959), .Y(n11962) );
  AOI22X1 U9014 ( .A(\lamb/scale_ls3/genblk1[1].mult/added[1] ), .B(n11964), 
        .C(n11143), .D(n11962), .Y(n11967) );
  AOI21X1 U9015 ( .A(n11967), .B(n11966), .C(n11965), .Y(n11978) );
  OAI21X1 U9016 ( .A(n10731), .B(\lamb/scale_bs3/genblk1[1].mult/added[3] ), 
        .C(\lamb/scale_bs3/genblk1[1].mult/added[1] ), .Y(n11969) );
  AOI21X1 U9017 ( .A(n11970), .B(n11969), .C(
        \lamb/scale_bs3/genblk1[1].mult/added[2] ), .Y(n11976) );
  INVX1 U9018 ( .A(n11971), .Y(n11972) );
  OAI21X1 U9019 ( .A(\lamb/scale_bs3/genblk1[1].mult/added[1] ), .B(n11973), 
        .C(n11972), .Y(n11975) );
  OAI21X1 U9020 ( .A(n11976), .B(n11975), .C(n11974), .Y(n11977) );
  HAX1 U9021 ( .A(n11978), .B(n11977), .YS(n13437) );
  INVX1 U9022 ( .A(n11979), .Y(n11980) );
  AOI22X1 U9023 ( .A(n11983), .B(n11982), .C(n11981), .D(n11980), .Y(n11986)
         );
  INVX1 U9024 ( .A(n11984), .Y(n11985) );
  NAND3X1 U9025 ( .A(n11987), .B(n11986), .C(n11985), .Y(n11988) );
  AOI22X1 U9026 ( .A(\lamb/scale_ls3/genblk1[0].mult/added[1] ), .B(n11991), 
        .C(\lamb/scale_ls3/genblk1[0].mult/added[2] ), .D(n10588), .Y(n11993)
         );
  NAND3X1 U9027 ( .A(n11994), .B(n11993), .C(n11992), .Y(n11996) );
  NAND2X1 U9028 ( .A(n11996), .B(n10677), .Y(n11997) );
  HAX1 U9029 ( .A(n10980), .B(n11997), .YS(n12061) );
  XNOR2X1 U9030 ( .A(n13437), .B(n12061), .Y(n12046) );
  HAX1 U9031 ( .A(n10843), .B(n12046), .YS(n12040) );
  OAI21X1 U9032 ( .A(n12080), .B(n12164), .C(n12040), .Y(n11999) );
  AOI21X1 U9033 ( .A(n12080), .B(n12164), .C(n11999), .Y(n12000) );
  INVX1 U9034 ( .A(n12000), .Y(n12001) );
  AOI21X1 U9035 ( .A(n13436), .B(n12101), .C(n12001), .Y(n12002) );
  OAI21X1 U9036 ( .A(n13436), .B(n12101), .C(n12002), .Y(n12003) );
  AOI21X1 U9037 ( .A(n12084), .B(n12144), .C(n12003), .Y(n12004) );
  OAI21X1 U9038 ( .A(n12084), .B(n12144), .C(n12004), .Y(n12822) );
  INVX1 U9039 ( .A(n12090), .Y(n12059) );
  HAX1 U9040 ( .A(n13458), .B(n12059), .YS(n12039) );
  INVX1 U9041 ( .A(n13436), .Y(n13439) );
  XNOR2X1 U9042 ( .A(n13439), .B(n10840), .Y(n12036) );
  INVX1 U9043 ( .A(n13437), .Y(n12010) );
  HAX1 U9044 ( .A(n12109), .B(n10842), .YS(n12034) );
  HAX1 U9045 ( .A(n12161), .B(n12132), .YS(n12060) );
  HAX1 U9046 ( .A(n13478), .B(n12060), .YS(n12026) );
  OAI21X1 U9047 ( .A(n12010), .B(n12034), .C(n12026), .Y(n12005) );
  AOI21X1 U9048 ( .A(n12010), .B(n12034), .C(n12005), .Y(n12006) );
  OAI21X1 U9049 ( .A(n12061), .B(n12036), .C(n10871), .Y(n12007) );
  AOI21X1 U9050 ( .A(n12061), .B(n12036), .C(n12007), .Y(n12008) );
  OAI21X1 U9051 ( .A(n10843), .B(n12039), .C(n12008), .Y(n12009) );
  AOI21X1 U9052 ( .A(n10843), .B(n12039), .C(n12009), .Y(n12800) );
  INVX1 U9053 ( .A(n10442), .Y(n13903) );
  HAX1 U9054 ( .A(n10842), .B(n12144), .YS(n12053) );
  INVX1 U9055 ( .A(n12053), .Y(n12112) );
  NAND2X1 U9056 ( .A(n13436), .B(n12010), .Y(n13430) );
  XNOR2X1 U9057 ( .A(n12109), .B(n13439), .Y(n12072) );
  HAX1 U9058 ( .A(n13458), .B(n10840), .YS(n12056) );
  HAX1 U9059 ( .A(n13437), .B(n13478), .YS(n13427) );
  XNOR2X1 U9060 ( .A(n13427), .B(n12132), .Y(n12105) );
  HAX1 U9061 ( .A(n13458), .B(n12010), .YS(n12117) );
  HAX1 U9062 ( .A(n12161), .B(n12117), .YS(n12108) );
  HAX1 U9063 ( .A(n13439), .B(n10843), .YS(n12153) );
  XNOR2X1 U9064 ( .A(n12108), .B(n12153), .Y(n12011) );
  INVX1 U9065 ( .A(n12061), .Y(n12113) );
  OR2X1 U9066 ( .A(n12011), .B(n12113), .Y(n12013) );
  NAND3X1 U9067 ( .A(n12105), .B(n12011), .C(n12113), .Y(n12012) );
  OAI21X1 U9068 ( .A(n12105), .B(n12013), .C(n12012), .Y(n12014) );
  OAI21X1 U9069 ( .A(n12072), .B(n12056), .C(n12014), .Y(n12015) );
  AOI21X1 U9070 ( .A(n12072), .B(n12056), .C(n12015), .Y(n12016) );
  OAI21X1 U9071 ( .A(n12112), .B(n10821), .C(n12016), .Y(n12017) );
  AOI21X1 U9072 ( .A(n12112), .B(n10821), .C(n12017), .Y(n12834) );
  INVX1 U9073 ( .A(n10450), .Y(n12431) );
  HAX1 U9074 ( .A(n10840), .B(n12080), .YS(n12150) );
  HAX1 U9075 ( .A(n13458), .B(n13439), .YS(n12098) );
  HAX1 U9076 ( .A(n10843), .B(n12161), .YS(n12125) );
  INVX1 U9077 ( .A(n12125), .Y(n12023) );
  INVX1 U9078 ( .A(n12045), .Y(n12057) );
  HAX1 U9079 ( .A(n10842), .B(n13427), .YS(n12018) );
  HAX1 U9080 ( .A(n12109), .B(n12061), .YS(n12151) );
  HAX1 U9081 ( .A(n12117), .B(n12151), .YS(n12127) );
  XNOR2X1 U9082 ( .A(n12127), .B(n12132), .Y(n12142) );
  AND2X1 U9083 ( .A(n12018), .B(n12142), .Y(n12020) );
  OAI21X1 U9084 ( .A(n12018), .B(n12142), .C(n12057), .Y(n12019) );
  OAI21X1 U9085 ( .A(n12057), .B(n12020), .C(n12019), .Y(n12021) );
  AOI21X1 U9086 ( .A(n12098), .B(n12023), .C(n12021), .Y(n12022) );
  OAI21X1 U9087 ( .A(n12098), .B(n12023), .C(n10867), .Y(n12024) );
  AOI21X1 U9088 ( .A(n12072), .B(n12150), .C(n12024), .Y(n12025) );
  OAI21X1 U9089 ( .A(n12072), .B(n12150), .C(n12025), .Y(n13586) );
  INVX1 U9090 ( .A(n10573), .Y(n12081) );
  HAX1 U9091 ( .A(n12072), .B(n12026), .YS(n12027) );
  OAI21X1 U9092 ( .A(n12127), .B(n12101), .C(n12027), .Y(n12028) );
  AOI21X1 U9093 ( .A(n12127), .B(n12101), .C(n12028), .Y(n12033) );
  HAX1 U9094 ( .A(n12046), .B(n12036), .YS(n12031) );
  HAX1 U9095 ( .A(n11196), .B(n12151), .YS(n12124) );
  HAX1 U9096 ( .A(n12124), .B(n12153), .YS(n12029) );
  MUX2X1 U9097 ( .B(n12031), .A(n12059), .S(n12029), .Y(n12030) );
  AOI21X1 U9098 ( .A(n12059), .B(n12031), .C(n12030), .Y(n12032) );
  HAX1 U9099 ( .A(n12035), .B(n12034), .YS(n12141) );
  HAX1 U9100 ( .A(n12061), .B(n12059), .YS(n12096) );
  HAX1 U9101 ( .A(n12161), .B(n12096), .YS(n12136) );
  FAX1 U9102 ( .A(n13429), .B(n12136), .C(n12036), .YS(n12042) );
  MUX2X1 U9103 ( .B(n12040), .A(n12039), .S(n12037), .Y(n12038) );
  AOI21X1 U9104 ( .A(n12040), .B(n12039), .C(n12038), .Y(n12041) );
  AOI21X1 U9105 ( .A(n10821), .B(n12141), .C(n10907), .Y(n12044) );
  OAI21X1 U9106 ( .A(n10821), .B(n12141), .C(n12044), .Y(n12853) );
  HAX1 U9107 ( .A(n12045), .B(n12153), .YS(n12147) );
  NAND2X1 U9108 ( .A(n12060), .B(n12046), .Y(n12050) );
  INVX1 U9109 ( .A(n12060), .Y(n12048) );
  INVX1 U9110 ( .A(n12046), .Y(n12047) );
  NAND3X1 U9111 ( .A(n12147), .B(n12048), .C(n12047), .Y(n12049) );
  OAI21X1 U9112 ( .A(n12147), .B(n12050), .C(n12049), .Y(n12051) );
  OAI21X1 U9113 ( .A(n12053), .B(n12072), .C(n12051), .Y(n12052) );
  AOI21X1 U9114 ( .A(n12053), .B(n12072), .C(n12052), .Y(n12054) );
  OAI21X1 U9115 ( .A(n12151), .B(n12056), .C(n10869), .Y(n12055) );
  AOI21X1 U9116 ( .A(n12151), .B(n12056), .C(n12055), .Y(n12850) );
  INVX1 U9117 ( .A(n10447), .Y(n12829) );
  HAX1 U9118 ( .A(n12109), .B(n10843), .YS(n12094) );
  HAX1 U9119 ( .A(n13427), .B(n12057), .YS(n12070) );
  HAX1 U9120 ( .A(n12059), .B(n10839), .YS(n12097) );
  INVX1 U9121 ( .A(n12097), .Y(n12067) );
  HAX1 U9122 ( .A(n13437), .B(n12060), .YS(n12064) );
  XNOR2X1 U9123 ( .A(n10842), .B(n12080), .Y(n12063) );
  HAX1 U9124 ( .A(n12061), .B(n12072), .YS(n12104) );
  MUX2X1 U9125 ( .B(n12063), .A(n12064), .S(n12104), .Y(n12062) );
  OAI21X1 U9126 ( .A(n12064), .B(n12063), .C(n12062), .Y(n12065) );
  AOI21X1 U9127 ( .A(n12127), .B(n12067), .C(n12065), .Y(n12066) );
  OAI21X1 U9128 ( .A(n12127), .B(n12067), .C(n10866), .Y(n12068) );
  AOI21X1 U9129 ( .A(n12094), .B(n12070), .C(n12068), .Y(n12069) );
  OAI21X1 U9130 ( .A(n12094), .B(n12070), .C(n12069), .Y(n12935) );
  INVX1 U9131 ( .A(n12935), .Y(n12809) );
  AOI21X1 U9132 ( .A(n10793), .B(n12810), .C(n12809), .Y(n13485) );
  HAX1 U9133 ( .A(n13439), .B(n12132), .YS(n12111) );
  XNOR2X1 U9134 ( .A(n13458), .B(n10842), .Y(n12082) );
  HAX1 U9135 ( .A(n12113), .B(n12082), .YS(n12160) );
  HAX1 U9136 ( .A(n13436), .B(n12160), .YS(n12077) );
  HAX1 U9137 ( .A(n10843), .B(n12072), .YS(n12074) );
  MUX2X1 U9138 ( .B(n13427), .A(n12084), .S(n12074), .Y(n12075) );
  AOI21X1 U9139 ( .A(n12084), .B(n13427), .C(n12075), .Y(n12076) );
  AOI21X1 U9140 ( .A(n12111), .B(n12080), .C(n10908), .Y(n12079) );
  OAI21X1 U9141 ( .A(n12111), .B(n12080), .C(n12079), .Y(n12771) );
  INVX1 U9142 ( .A(n12771), .Y(n12833) );
  AOI21X1 U9143 ( .A(n12081), .B(n10691), .C(n13483), .Y(n12925) );
  INVX1 U9144 ( .A(n12098), .Y(n13426) );
  HAX1 U9145 ( .A(n13426), .B(n12132), .YS(n12091) );
  NAND2X1 U9146 ( .A(n12091), .B(n12090), .Y(n12088) );
  INVX1 U9147 ( .A(n12151), .Y(n12154) );
  HAX1 U9148 ( .A(n12154), .B(n12082), .YS(n12139) );
  INVX1 U9149 ( .A(n12084), .Y(n12121) );
  XNOR2X1 U9150 ( .A(n13478), .B(n12121), .Y(n12128) );
  HAX1 U9151 ( .A(n12113), .B(n12128), .YS(n12085) );
  MUX2X1 U9152 ( .B(n12083), .A(n12139), .S(n12085), .Y(n12086) );
  AOI21X1 U9153 ( .A(n12139), .B(n12083), .C(n12086), .Y(n12087) );
  NAND2X1 U9154 ( .A(n12088), .B(n10880), .Y(n12093) );
  HAX1 U9155 ( .A(n13426), .B(n13427), .YS(n12110) );
  HAX1 U9156 ( .A(n12110), .B(n12094), .YS(n12089) );
  MUX2X1 U9157 ( .B(n12091), .A(n12090), .S(n12089), .Y(n12092) );
  OR2X1 U9158 ( .A(n12093), .B(n12092), .Y(n12964) );
  INVX1 U9159 ( .A(n12094), .Y(n12095) );
  HAX1 U9160 ( .A(n13478), .B(n12095), .YS(n12135) );
  HAX1 U9161 ( .A(n13437), .B(n12097), .YS(n12155) );
  FAX1 U9162 ( .A(n12109), .B(n12098), .C(n12155), .YS(n12099) );
  AOI21X1 U9163 ( .A(n12126), .B(n12101), .C(n12099), .Y(n12100) );
  OAI21X1 U9164 ( .A(n12126), .B(n12101), .C(n10870), .Y(n12102) );
  AOI21X1 U9165 ( .A(n12105), .B(n12104), .C(n12102), .Y(n12103) );
  OAI21X1 U9166 ( .A(n12105), .B(n12104), .C(n12103), .Y(n12106) );
  AOI21X1 U9167 ( .A(n12135), .B(n12108), .C(n12106), .Y(n12107) );
  OAI21X1 U9168 ( .A(n12135), .B(n12108), .C(n12107), .Y(n13896) );
  INVX1 U9169 ( .A(n13896), .Y(n13891) );
  AOI21X1 U9170 ( .A(n11060), .B(n12964), .C(n13891), .Y(n12927) );
  XNOR2X1 U9171 ( .A(n12110), .B(n12109), .Y(n12120) );
  HAX1 U9172 ( .A(n12111), .B(n12136), .YS(n12116) );
  HAX1 U9173 ( .A(n12113), .B(n12112), .YS(n12114) );
  MUX2X1 U9174 ( .B(n12116), .A(n12117), .S(n12114), .Y(n12115) );
  OAI21X1 U9175 ( .A(n12117), .B(n12116), .C(n12115), .Y(n12118) );
  AOI21X1 U9176 ( .A(n12121), .B(n12120), .C(n12118), .Y(n12119) );
  OAI21X1 U9177 ( .A(n12121), .B(n12120), .C(n10868), .Y(n12122) );
  AOI21X1 U9178 ( .A(n12125), .B(n12124), .C(n12122), .Y(n12123) );
  OAI21X1 U9179 ( .A(n12125), .B(n12124), .C(n12123), .Y(n13488) );
  INVX1 U9180 ( .A(n12126), .Y(n12131) );
  HAX1 U9181 ( .A(n12128), .B(n12127), .YS(n12129) );
  AOI21X1 U9182 ( .A(n12132), .B(n12131), .C(n12129), .Y(n12130) );
  OAI21X1 U9183 ( .A(n12132), .B(n12131), .C(n12130), .Y(n12133) );
  AOI21X1 U9184 ( .A(n12136), .B(n12135), .C(n12133), .Y(n12134) );
  OAI21X1 U9185 ( .A(n12136), .B(n12135), .C(n12134), .Y(n12137) );
  AOI21X1 U9186 ( .A(n12144), .B(n12139), .C(n12137), .Y(n12138) );
  OAI21X1 U9187 ( .A(n12144), .B(n12139), .C(n12138), .Y(n12803) );
  INVX1 U9188 ( .A(n12803), .Y(n13487) );
  AOI21X1 U9189 ( .A(n10404), .B(n13488), .C(n13487), .Y(n12140) );
  INVX1 U9190 ( .A(n12140), .Y(n12152) );
  INVX1 U9191 ( .A(n12141), .Y(n12145) );
  MUX2X1 U9192 ( .B(n12144), .A(n12145), .S(n12142), .Y(n12143) );
  AOI21X1 U9193 ( .A(n12145), .B(n12144), .C(n12143), .Y(n12146) );
  AOI21X1 U9194 ( .A(n12151), .B(n12150), .C(n10906), .Y(n12149) );
  OAI21X1 U9195 ( .A(n12151), .B(n12150), .C(n12149), .Y(n12804) );
  NAND2X1 U9196 ( .A(n13695), .B(n10582), .Y(n12772) );
  INVX1 U9197 ( .A(n12772), .Y(n12165) );
  INVX1 U9198 ( .A(n10437), .Y(n12795) );
  INVX1 U9199 ( .A(n10570), .Y(n13893) );
  HAX1 U9200 ( .A(n12154), .B(n12153), .YS(n12157) );
  OAI21X1 U9201 ( .A(n13429), .B(n12157), .C(n12155), .Y(n12156) );
  AOI21X1 U9202 ( .A(n13429), .B(n12157), .C(n12156), .Y(n12158) );
  OAI21X1 U9203 ( .A(n12161), .B(n12160), .C(n12158), .Y(n12159) );
  AOI21X1 U9204 ( .A(n12161), .B(n12160), .C(n12159), .Y(n12162) );
  OAI21X1 U9205 ( .A(n13436), .B(n12164), .C(n12162), .Y(n12163) );
  AOI21X1 U9206 ( .A(n13436), .B(n12164), .C(n12163), .Y(n12849) );
  INVX1 U9207 ( .A(n12856), .Y(n12936) );
  OAI21X1 U9208 ( .A(n12809), .B(n12936), .C(n12827), .Y(n12938) );
  NAND2X1 U9209 ( .A(n13896), .B(n12938), .Y(n12943) );
  NAND2X1 U9210 ( .A(n13893), .B(n12943), .Y(n12950) );
  AND2X1 U9211 ( .A(n12165), .B(n12950), .Y(\forney/m0/logA [3]) );
  INVX1 U9212 ( .A(n12964), .Y(n13486) );
  AOI21X1 U9213 ( .A(n12771), .B(n10409), .C(n10450), .Y(n12812) );
  OAI21X1 U9214 ( .A(n13486), .B(n12812), .C(n13896), .Y(n12821) );
  OAI21X1 U9215 ( .A(n11172), .B(n12821), .C(n13695), .Y(n13001) );
  INVX1 U9216 ( .A(n10564), .Y(n13602) );
  INVX1 U9217 ( .A(n10546), .Y(n12832) );
  NAND2X1 U9218 ( .A(n11161), .B(n12829), .Y(n12166) );
  AOI21X1 U9219 ( .A(n12832), .B(n12166), .C(n10573), .Y(n12167) );
  INVX1 U9220 ( .A(n12853), .Y(n12807) );
  AOI21X1 U9221 ( .A(n12167), .B(n11079), .C(n13483), .Y(n12837) );
  NOR2X1 U9222 ( .A(n10793), .B(n12809), .Y(n12963) );
  NAND2X1 U9223 ( .A(n12963), .B(n13586), .Y(n12852) );
  NAND2X1 U9224 ( .A(n12964), .B(n10986), .Y(n12966) );
  NAND2X1 U9225 ( .A(n13896), .B(n12966), .Y(n12968) );
  NAND2X1 U9226 ( .A(n13488), .B(n12968), .Y(n12971) );
  NAND2X1 U9227 ( .A(n13602), .B(n12971), .Y(n12974) );
  NAND2X1 U9228 ( .A(n11164), .B(n12997), .Y(n12630) );
  INVX1 U9229 ( .A(n13001), .Y(n12993) );
  NAND2X1 U9230 ( .A(n12993), .B(n12997), .Y(n12631) );
  NAND3X1 U9231 ( .A(n12771), .B(n13586), .C(n11079), .Y(n12790) );
  NAND2X1 U9232 ( .A(n12431), .B(n12790), .Y(n12793) );
  AOI21X1 U9233 ( .A(n12964), .B(n12793), .C(n13891), .Y(n12169) );
  INVX1 U9234 ( .A(n12169), .Y(n12797) );
  INVX1 U9235 ( .A(n10576), .Y(n12998) );
  AOI21X1 U9236 ( .A(n13003), .B(n12631), .C(n12998), .Y(n12994) );
  NOR3X1 U9237 ( .A(\lamb/scale_ds3/genblk1[2].mult/added[3] ), .B(
        \add_x_121/n1 ), .C(\lamb/scale_ds3/genblk1[2].mult/added[4] ), .Y(
        n12398) );
  INVX1 U9238 ( .A(\lamb/scale_ds3/genblk1[2].mult/added[3] ), .Y(n12170) );
  NOR2X1 U9239 ( .A(\add_x_121/n1 ), .B(
        \lamb/scale_ds3/genblk1[2].mult/added[4] ), .Y(n12380) );
  OR2X1 U9240 ( .A(n12170), .B(n12380), .Y(n12400) );
  NOR2X1 U9241 ( .A(\lamb/scale_ds3/genblk1[2].mult/added[1] ), .B(n12400), 
        .Y(n12179) );
  NAND2X1 U9242 ( .A(n12179), .B(n11098), .Y(n12415) );
  NAND2X1 U9243 ( .A(\lamb/scale_ds3/genblk1[2].mult/added[2] ), .B(n12415), 
        .Y(n12175) );
  INVX1 U9244 ( .A(\lamb/scale_ds3/genblk1[2].mult/added[2] ), .Y(n12173) );
  NAND3X1 U9245 ( .A(\lamb/scale_ds3/genblk1[2].mult/added[3] ), .B(
        \add_x_121/n1 ), .C(\lamb/scale_ds3/genblk1[2].mult/added[4] ), .Y(
        n12176) );
  NAND2X1 U9246 ( .A(n12170), .B(n11098), .Y(n12171) );
  NAND2X1 U9247 ( .A(n12417), .B(\lamb/scale_ds3/genblk1[2].mult/added[1] ), 
        .Y(n12172) );
  NAND3X1 U9248 ( .A(n12173), .B(n12176), .C(n12172), .Y(n12174) );
  OAI21X1 U9249 ( .A(n12398), .B(n12175), .C(n12174), .Y(n12383) );
  NAND2X1 U9250 ( .A(\lamb/scale_ds3/genblk1[2].mult/added[1] ), .B(
        \lamb/scale_ds3/genblk1[2].mult/added[2] ), .Y(n12397) );
  INVX1 U9251 ( .A(n12397), .Y(n12177) );
  AOI21X1 U9252 ( .A(n12177), .B(n12176), .C(n12398), .Y(n12381) );
  NAND3X1 U9253 ( .A(n12178), .B(n12179), .C(
        \lamb/scale_ds3/genblk1[2].mult/added[2] ), .Y(n12402) );
  NAND3X1 U9254 ( .A(n12383), .B(n11018), .C(n10433), .Y(n12283) );
  NAND3X1 U9255 ( .A(\lamb/scale_ts2/genblk1[1].mult/added[3] ), .B(
        \add_x_131/n1 ), .C(\lamb/scale_ts2/genblk1[1].mult/added[4] ), .Y(
        n12243) );
  NOR3X1 U9256 ( .A(\lamb/scale_ts2/genblk1[1].mult/added[3] ), .B(
        \add_x_131/n1 ), .C(\lamb/scale_ts2/genblk1[1].mult/added[4] ), .Y(
        n12181) );
  AOI21X1 U9257 ( .A(\lamb/scale_ts2/genblk1[1].mult/added[2] ), .B(n10519), 
        .C(n12181), .Y(n12180) );
  INVX1 U9258 ( .A(\lamb/scale_ts2/genblk1[1].mult/added[3] ), .Y(n12240) );
  NAND2X1 U9259 ( .A(\add_x_131/n1 ), .B(
        \lamb/scale_ts2/genblk1[1].mult/added[4] ), .Y(n12237) );
  OAI21X1 U9260 ( .A(\add_x_131/n1 ), .B(
        \lamb/scale_ts2/genblk1[1].mult/added[4] ), .C(n12237), .Y(n12242) );
  INVX1 U9261 ( .A(n12242), .Y(n12256) );
  INVX1 U9262 ( .A(\lamb/scale_ts2/genblk1[1].mult/added[1] ), .Y(n12182) );
  AOI22X1 U9263 ( .A(\lamb/scale_ts2/genblk1[1].mult/added[1] ), .B(n12180), 
        .C(n12264), .D(n12182), .Y(n12216) );
  INVX1 U9264 ( .A(n10519), .Y(n12184) );
  INVX1 U9265 ( .A(n12181), .Y(n12266) );
  NAND3X1 U9266 ( .A(n12256), .B(\lamb/scale_ts2/genblk1[1].mult/added[3] ), 
        .C(n12182), .Y(n12271) );
  NAND3X1 U9267 ( .A(n12266), .B(n12271), .C(
        \lamb/scale_ts2/genblk1[1].mult/added[2] ), .Y(n12183) );
  OAI21X1 U9268 ( .A(\lamb/scale_ts2/genblk1[1].mult/added[2] ), .B(n12184), 
        .C(n12183), .Y(n12265) );
  INVX1 U9269 ( .A(n12659), .Y(n12663) );
  AOI22X1 U9270 ( .A(n10851), .B(n13367), .C(n12663), .D(n12682), .Y(n13284)
         );
  NOR3X1 U9271 ( .A(\lamb/scale_ts0/genblk1[0].mult/added[4] ), .B(
        \add_x_154/n1 ), .C(\lamb/scale_ts0/genblk1[0].mult/added[3] ), .Y(
        n12198) );
  NAND3X1 U9272 ( .A(\lamb/scale_ts0/genblk1[0].mult/added[4] ), .B(
        \add_x_154/n1 ), .C(\lamb/scale_ts0/genblk1[0].mult/added[3] ), .Y(
        n12185) );
  OAI21X1 U9273 ( .A(n12201), .B(n12198), .C(n12185), .Y(n12192) );
  INVX1 U9274 ( .A(n12185), .Y(n12194) );
  INVX1 U9275 ( .A(\lamb/scale_ts0/genblk1[0].mult/added[2] ), .Y(n12203) );
  AOI22X1 U9276 ( .A(\lamb/scale_ts0/genblk1[0].mult/added[2] ), .B(n12198), 
        .C(n12194), .D(n12203), .Y(n12188) );
  AOI21X1 U9277 ( .A(\add_x_154/n1 ), .B(
        \lamb/scale_ts0/genblk1[0].mult/added[4] ), .C(
        \lamb/scale_ts0/genblk1[0].mult/added[3] ), .Y(n12191) );
  OR2X1 U9278 ( .A(\lamb/scale_ts0/genblk1[0].mult/added[4] ), .B(
        \add_x_154/n1 ), .Y(n12186) );
  AND2X1 U9279 ( .A(n12191), .B(n12186), .Y(n12211) );
  NAND2X1 U9280 ( .A(n12211), .B(n10702), .Y(n12197) );
  AND2X1 U9281 ( .A(\lamb/scale_ts0/genblk1[0].mult/added[4] ), .B(
        \add_x_154/n1 ), .Y(n12187) );
  NOR3X1 U9282 ( .A(\lamb/scale_ts0/genblk1[0].mult/added[1] ), .B(n12187), 
        .C(n11184), .Y(n12212) );
  NAND2X1 U9283 ( .A(\lamb/scale_ts0/genblk1[0].mult/added[2] ), .B(n12212), 
        .Y(n12195) );
  NAND3X1 U9284 ( .A(n12188), .B(n12197), .C(n12195), .Y(n12189) );
  AOI21X1 U9285 ( .A(\lamb/scale_ts0/genblk1[0].mult/added[1] ), .B(n12192), 
        .C(n12189), .Y(n13356) );
  INVX1 U9286 ( .A(n11119), .Y(n13355) );
  NAND2X1 U9287 ( .A(n12659), .B(n12664), .Y(n12190) );
  AOI21X1 U9288 ( .A(n12665), .B(n12190), .C(n12667), .Y(n12673) );
  AOI21X1 U9289 ( .A(n12659), .B(n11133), .C(n12664), .Y(n12672) );
  INVX1 U9290 ( .A(n10465), .Y(n12335) );
  AND2X1 U9291 ( .A(n13355), .B(n12335), .Y(n12724) );
  AOI22X1 U9292 ( .A(n10795), .B(n13235), .C(n12724), .D(n13224), .Y(n13187)
         );
  AOI22X1 U9293 ( .A(n10851), .B(n12293), .C(n12667), .D(n12682), .Y(n13280)
         );
  INVX1 U9294 ( .A(\lamb/scale_ts0/genblk1[0].mult/added[1] ), .Y(n12205) );
  INVX1 U9295 ( .A(n12191), .Y(n12206) );
  OAI21X1 U9296 ( .A(n12205), .B(n10663), .C(n12192), .Y(n12193) );
  NAND2X1 U9297 ( .A(n12194), .B(n10702), .Y(n12196) );
  NAND2X1 U9298 ( .A(n12335), .B(n13924), .Y(n13359) );
  AOI22X1 U9299 ( .A(n10851), .B(n13370), .C(n12665), .D(n12682), .Y(n13288)
         );
  NAND2X1 U9300 ( .A(n12197), .B(n12196), .Y(n12202) );
  INVX1 U9301 ( .A(n12198), .Y(n12199) );
  OAI21X1 U9302 ( .A(n12199), .B(n12205), .C(n10663), .Y(n12200) );
  AOI22X1 U9303 ( .A(\lamb/scale_ts0/genblk1[0].mult/added[2] ), .B(n12202), 
        .C(n10702), .D(n12200), .Y(n13354) );
  AOI22X1 U9304 ( .A(n12205), .B(n10663), .C(n12203), .D(n11184), .Y(n12207)
         );
  NAND2X1 U9305 ( .A(n12206), .B(n12201), .Y(n12208) );
  NAND2X1 U9306 ( .A(n12207), .B(n12208), .Y(n13927) );
  NOR2X1 U9307 ( .A(n10800), .B(n10805), .Y(n13179) );
  AOI22X1 U9308 ( .A(n10851), .B(n13826), .C(n12670), .D(n12682), .Y(n13289)
         );
  INVX1 U9309 ( .A(n12208), .Y(n12210) );
  AOI22X1 U9310 ( .A(\lamb/scale_ts0/genblk1[0].mult/added[1] ), .B(n12211), 
        .C(n12210), .D(n11184), .Y(n12213) );
  INVX1 U9311 ( .A(n10474), .Y(n12725) );
  AOI22X1 U9312 ( .A(n13235), .B(n10797), .C(n12725), .D(n10809), .Y(n13946)
         );
  NAND3X1 U9313 ( .A(n10703), .B(n13179), .C(n10832), .Y(n12214) );
  AOI21X1 U9314 ( .A(n12216), .B(n12265), .C(n11116), .Y(n12225) );
  NAND3X1 U9315 ( .A(\lamb/scale_ds2/genblk1[1].mult/added[2] ), .B(
        \lamb/scale_ds2/genblk1[1].mult/added[3] ), .C(n12217), .Y(n12232) );
  AOI21X1 U9316 ( .A(\lamb/scale_ds2/genblk1[1].mult/added[3] ), .B(n12217), 
        .C(\lamb/scale_ds2/genblk1[1].mult/added[2] ), .Y(n12219) );
  OR2X1 U9317 ( .A(\add_x_135/n1 ), .B(
        \lamb/scale_ds2/genblk1[1].mult/added[4] ), .Y(n12228) );
  OR2X1 U9318 ( .A(n12228), .B(\lamb/scale_ds2/genblk1[1].mult/added[3] ), .Y(
        n12221) );
  NAND2X1 U9319 ( .A(n12232), .B(n11016), .Y(n12218) );
  INVX1 U9320 ( .A(\lamb/scale_ds2/genblk1[1].mult/added[1] ), .Y(n12233) );
  NAND2X1 U9321 ( .A(n10988), .B(n12228), .Y(n12275) );
  INVX1 U9322 ( .A(n12275), .Y(n12230) );
  AND2X1 U9323 ( .A(n12233), .B(n12230), .Y(n12220) );
  INVX1 U9324 ( .A(\lamb/scale_ds2/genblk1[1].mult/added[3] ), .Y(n12227) );
  AOI22X1 U9325 ( .A(\lamb/scale_ds2/genblk1[1].mult/added[1] ), .B(n12218), 
        .C(n12220), .D(n12227), .Y(n12223) );
  INVX1 U9326 ( .A(n12219), .Y(n12222) );
  NAND2X1 U9327 ( .A(\lamb/scale_ds2/genblk1[1].mult/added[3] ), .B(n12220), 
        .Y(n12279) );
  NAND3X1 U9328 ( .A(\lamb/scale_ds2/genblk1[1].mult/added[2] ), .B(n12279), 
        .C(n12221), .Y(n12254) );
  AOI21X1 U9329 ( .A(n12223), .B(n10652), .C(n11209), .Y(n12224) );
  NAND2X1 U9330 ( .A(\lamb/scale_ds2/genblk1[1].mult/added[2] ), .B(
        \lamb/scale_ds2/genblk1[1].mult/added[3] ), .Y(n12273) );
  NAND3X1 U9331 ( .A(\add_x_135/n1 ), .B(
        \lamb/scale_ds2/genblk1[1].mult/added[4] ), .C(n12227), .Y(n12226) );
  OAI21X1 U9332 ( .A(n12228), .B(n12227), .C(n12226), .Y(n12278) );
  AOI21X1 U9333 ( .A(\lamb/scale_ds2/genblk1[1].mult/added[1] ), .B(n10924), 
        .C(n12278), .Y(n12231) );
  OAI21X1 U9334 ( .A(\lamb/scale_ds2/genblk1[1].mult/added[2] ), .B(n12231), 
        .C(n11021), .Y(n12236) );
  NAND2X1 U9335 ( .A(n12233), .B(n12232), .Y(n12252) );
  INVX1 U9336 ( .A(n12252), .Y(n12234) );
  INVX1 U9337 ( .A(n12278), .Y(n12250) );
  AOI22X1 U9338 ( .A(\lamb/scale_ds2/genblk1[1].mult/added[1] ), .B(n10652), 
        .C(n12234), .D(n12250), .Y(n12235) );
  AOI21X1 U9339 ( .A(n12273), .B(n12236), .C(n12235), .Y(n12248) );
  INVX1 U9340 ( .A(n12237), .Y(n12239) );
  NOR2X1 U9341 ( .A(n12240), .B(\lamb/scale_ts2/genblk1[1].mult/added[1] ), 
        .Y(n12238) );
  NAND3X1 U9342 ( .A(\lamb/scale_ts2/genblk1[1].mult/added[2] ), .B(n12239), 
        .C(n12238), .Y(n12259) );
  OR2X1 U9343 ( .A(n12242), .B(\lamb/scale_ts2/genblk1[1].mult/added[2] ), .Y(
        n12263) );
  AND2X1 U9344 ( .A(n12266), .B(n12265), .Y(n12257) );
  OAI21X1 U9345 ( .A(n12240), .B(n12263), .C(n12257), .Y(n12241) );
  AOI22X1 U9346 ( .A(\lamb/scale_ts2/genblk1[1].mult/added[2] ), .B(n12264), 
        .C(\lamb/scale_ts2/genblk1[1].mult/added[1] ), .D(n12241), .Y(n12245)
         );
  NAND2X1 U9347 ( .A(\lamb/scale_ts2/genblk1[1].mult/added[2] ), .B(
        \lamb/scale_ts2/genblk1[1].mult/added[1] ), .Y(n12255) );
  NAND3X1 U9348 ( .A(n12259), .B(n12245), .C(n12244), .Y(n12246) );
  NAND2X1 U9349 ( .A(n12270), .B(n12246), .Y(n12247) );
  OAI21X1 U9350 ( .A(n12248), .B(n11209), .C(n12247), .Y(n13077) );
  NAND3X1 U9351 ( .A(n12250), .B(\lamb/scale_ds2/genblk1[1].mult/added[1] ), 
        .C(n11021), .Y(n12251) );
  AOI22X1 U9352 ( .A(n12254), .B(n11016), .C(n12252), .D(n12251), .Y(n12262)
         );
  AOI22X1 U9353 ( .A(n12256), .B(n10960), .C(
        \lamb/scale_ts2/genblk1[1].mult/added[1] ), .D(n12267), .Y(n12258) );
  NAND2X1 U9354 ( .A(n12270), .B(n12260), .Y(n12261) );
  OAI21X1 U9355 ( .A(n12262), .B(n11209), .C(n12261), .Y(n13072) );
  NAND3X1 U9356 ( .A(n12265), .B(n11000), .C(n12263), .Y(n12269) );
  AND2X1 U9357 ( .A(\lamb/scale_ts2/genblk1[1].mult/added[2] ), .B(n12266), 
        .Y(n12268) );
  AOI22X1 U9358 ( .A(\lamb/scale_ts2/genblk1[1].mult/added[1] ), .B(n12269), 
        .C(n12268), .D(n12267), .Y(n12272) );
  AOI21X1 U9359 ( .A(n12272), .B(n12271), .C(n11116), .Y(n12282) );
  INVX1 U9360 ( .A(n12273), .Y(n12276) );
  OAI21X1 U9361 ( .A(n12276), .B(n12275), .C(n10652), .Y(n12277) );
  AOI22X1 U9362 ( .A(\lamb/scale_ds2/genblk1[1].mult/added[2] ), .B(n12278), 
        .C(\lamb/scale_ds2/genblk1[1].mult/added[1] ), .D(n12277), .Y(n12280)
         );
  AOI21X1 U9363 ( .A(n12280), .B(n12279), .C(n11209), .Y(n12281) );
  AOI21X1 U9364 ( .A(n13070), .B(n10650), .C(n13081), .Y(n13067) );
  NAND2X1 U9365 ( .A(n10724), .B(n13072), .Y(n13065) );
  INVX1 U9366 ( .A(n13065), .Y(n13078) );
  NOR2X1 U9367 ( .A(n13077), .B(n13078), .Y(n13076) );
  NAND2X1 U9368 ( .A(n12283), .B(n11155), .Y(n12374) );
  INVX1 U9369 ( .A(\lamb/scale_ts3/genblk1[2].mult/added[3] ), .Y(n12288) );
  AOI22X1 U9370 ( .A(n12289), .B(\lamb/scale_ts3/genblk1[2].mult/added[3] ), 
        .C(n11182), .D(n10428), .Y(n12376) );
  NOR2X1 U9371 ( .A(\lamb/scale_ts3/genblk1[2].mult/added[1] ), .B(n12391), 
        .Y(n12285) );
  NAND2X1 U9372 ( .A(\lamb/scale_ts3/genblk1[2].mult/added[2] ), .B(n11182), 
        .Y(n12392) );
  INVX1 U9373 ( .A(n12392), .Y(n12284) );
  NOR2X1 U9374 ( .A(n10682), .B(n12288), .Y(n12287) );
  NAND2X1 U9375 ( .A(n12285), .B(n10682), .Y(n12408) );
  NAND3X1 U9376 ( .A(\lamb/scale_ts3/genblk1[2].mult/added[2] ), .B(n12408), 
        .C(n11182), .Y(n12286) );
  OAI21X1 U9377 ( .A(\lamb/scale_ts3/genblk1[2].mult/added[2] ), .B(n12287), 
        .C(n12286), .Y(n12379) );
  NAND2X1 U9378 ( .A(n10682), .B(n12288), .Y(n12290) );
  INVX1 U9379 ( .A(\lamb/scale_ts3/genblk1[2].mult/added[1] ), .Y(n12386) );
  OR2X1 U9380 ( .A(n10516), .B(n12386), .Y(n12291) );
  NAND3X1 U9381 ( .A(n12394), .B(n12379), .C(n12291), .Y(n12372) );
  AOI22X1 U9382 ( .A(n12293), .B(n11713), .C(n12292), .D(n10809), .Y(n12689)
         );
  NOR3X1 U9383 ( .A(\add_x_144/n1 ), .B(
        \lamb/scale_ts1/genblk1[1].mult/added[4] ), .C(
        \lamb/scale_ts1/genblk1[1].mult/added[3] ), .Y(n12319) );
  AOI21X1 U9384 ( .A(\lamb/scale_ts1/genblk1[1].mult/added[4] ), .B(
        \add_x_144/n1 ), .C(\lamb/scale_ts1/genblk1[1].mult/added[3] ), .Y(
        n12295) );
  OR2X1 U9385 ( .A(\add_x_144/n1 ), .B(
        \lamb/scale_ts1/genblk1[1].mult/added[4] ), .Y(n12296) );
  AND2X1 U9386 ( .A(n12295), .B(n12296), .Y(n12353) );
  NAND2X1 U9387 ( .A(\lamb/scale_ts1/genblk1[1].mult/added[1] ), .B(
        \lamb/scale_ts1/genblk1[1].mult/added[2] ), .Y(n12322) );
  INVX1 U9388 ( .A(n12322), .Y(n12294) );
  NAND3X1 U9389 ( .A(\add_x_144/n1 ), .B(
        \lamb/scale_ts1/genblk1[1].mult/added[4] ), .C(
        \lamb/scale_ts1/genblk1[1].mult/added[3] ), .Y(n12301) );
  OAI21X1 U9390 ( .A(\lamb/scale_ts1/genblk1[1].mult/added[1] ), .B(n12353), 
        .C(n11022), .Y(n12345) );
  INVX1 U9391 ( .A(n12345), .Y(n12300) );
  INVX1 U9392 ( .A(n12295), .Y(n12321) );
  AND2X1 U9393 ( .A(n12321), .B(n10653), .Y(n12354) );
  INVX1 U9394 ( .A(\lamb/scale_ts1/genblk1[1].mult/added[2] ), .Y(n12350) );
  NOR2X1 U9395 ( .A(n12350), .B(n12319), .Y(n12349) );
  OR2X1 U9396 ( .A(\lamb/scale_ts1/genblk1[1].mult/added[1] ), .B(n10653), .Y(
        n12320) );
  INVX1 U9397 ( .A(n12320), .Y(n12298) );
  NAND2X1 U9398 ( .A(\add_x_144/n1 ), .B(
        \lamb/scale_ts1/genblk1[1].mult/added[4] ), .Y(n12297) );
  AOI22X1 U9399 ( .A(n12349), .B(n11057), .C(n10618), .D(n12350), .Y(n12299)
         );
  AOI21X1 U9400 ( .A(n12300), .B(n12354), .C(n12299), .Y(n12344) );
  NOR2X1 U9401 ( .A(\lamb/scale_ts1/genblk1[1].mult/added[1] ), .B(n10618), 
        .Y(n12318) );
  INVX1 U9402 ( .A(n12318), .Y(n12303) );
  NAND3X1 U9403 ( .A(n12344), .B(n12303), .C(n11022), .Y(n12306) );
  AOI21X1 U9404 ( .A(n10795), .B(n10657), .C(n10797), .Y(n13282) );
  INVX1 U9405 ( .A(n12304), .Y(n12305) );
  AOI21X1 U9406 ( .A(n10424), .B(n10430), .C(n12305), .Y(n12356) );
  OAI21X1 U9407 ( .A(n12319), .B(n12306), .C(n11147), .Y(n12317) );
  NAND3X1 U9408 ( .A(\lamb/scale_ds1/genblk1[1].mult/added[3] ), .B(
        \add_x_148/n1 ), .C(\lamb/scale_ds1/genblk1[1].mult/added[4] ), .Y(
        n12308) );
  NOR3X1 U9409 ( .A(\lamb/scale_ds1/genblk1[1].mult/added[3] ), .B(
        \add_x_148/n1 ), .C(\lamb/scale_ds1/genblk1[1].mult/added[4] ), .Y(
        n12307) );
  AOI21X1 U9410 ( .A(n12339), .B(n12308), .C(n12307), .Y(n12340) );
  INVX1 U9411 ( .A(\lamb/scale_ds1/genblk1[1].mult/added[3] ), .Y(n12329) );
  INVX1 U9412 ( .A(n12307), .Y(n12311) );
  OR2X1 U9413 ( .A(\add_x_148/n1 ), .B(
        \lamb/scale_ds1/genblk1[1].mult/added[4] ), .Y(n12328) );
  NAND2X1 U9414 ( .A(n12311), .B(n10987), .Y(n12326) );
  AOI21X1 U9415 ( .A(n12329), .B(n11183), .C(n12326), .Y(n12360) );
  INVX1 U9416 ( .A(n12308), .Y(n12312) );
  INVX1 U9417 ( .A(\lamb/scale_ds1/genblk1[1].mult/added[1] ), .Y(n12309) );
  AOI22X1 U9418 ( .A(\lamb/scale_ds1/genblk1[1].mult/added[1] ), .B(n10631), 
        .C(n12312), .D(n12309), .Y(n12314) );
  NAND3X1 U9419 ( .A(n11183), .B(n10754), .C(n12310), .Y(n12367) );
  INVX1 U9420 ( .A(n12367), .Y(n12313) );
  NAND2X1 U9421 ( .A(\lamb/scale_ds1/genblk1[1].mult/added[2] ), .B(n12311), 
        .Y(n12327) );
  OR2X1 U9422 ( .A(n12312), .B(\lamb/scale_ds1/genblk1[1].mult/added[2] ), .Y(
        n12364) );
  OAI21X1 U9423 ( .A(n12313), .B(n12327), .C(n12364), .Y(n12341) );
  NAND3X1 U9424 ( .A(n11053), .B(n12314), .C(n12341), .Y(n12315) );
  NAND2X1 U9425 ( .A(n12315), .B(n12335), .Y(n12316) );
  HAX1 U9426 ( .A(n12317), .B(n12316), .YS(n13933) );
  INVX1 U9427 ( .A(n13933), .Y(n13206) );
  AOI22X1 U9428 ( .A(n11227), .B(n10444), .C(n13206), .D(n13841), .Y(n13046)
         );
  AOI22X1 U9429 ( .A(n13235), .B(n13269), .C(n13342), .D(n10809), .Y(n13175)
         );
  OAI21X1 U9430 ( .A(n12318), .B(n12353), .C(
        \lamb/scale_ts1/genblk1[1].mult/added[2] ), .Y(n12324) );
  NAND3X1 U9431 ( .A(n12322), .B(n12321), .C(n12320), .Y(n12323) );
  NAND3X1 U9432 ( .A(n12324), .B(n10999), .C(n12323), .Y(n12325) );
  NAND2X1 U9433 ( .A(n11147), .B(n12325), .Y(n12337) );
  INVX1 U9434 ( .A(n12326), .Y(n12333) );
  NAND2X1 U9435 ( .A(\lamb/scale_ds1/genblk1[1].mult/added[1] ), .B(n12327), 
        .Y(n12361) );
  NAND3X1 U9436 ( .A(n12329), .B(n12328), .C(n11183), .Y(n12338) );
  OAI21X1 U9437 ( .A(\lamb/scale_ds1/genblk1[1].mult/added[1] ), .B(n11183), 
        .C(n12338), .Y(n12331) );
  AOI22X1 U9438 ( .A(\lamb/scale_ds1/genblk1[1].mult/added[2] ), .B(n12331), 
        .C(n10631), .D(n10754), .Y(n12332) );
  OAI21X1 U9439 ( .A(n12333), .B(n12361), .C(n12332), .Y(n12334) );
  HAX1 U9440 ( .A(n12337), .B(n10973), .YS(n13937) );
  INVX1 U9441 ( .A(n13937), .Y(n13204) );
  AOI22X1 U9442 ( .A(n11227), .B(n10726), .C(n13204), .D(n13841), .Y(n13038)
         );
  INVX1 U9443 ( .A(n13038), .Y(n13044) );
  AND2X1 U9444 ( .A(n10829), .B(n13044), .Y(n13037) );
  INVX1 U9445 ( .A(n13267), .Y(n13272) );
  AOI22X1 U9446 ( .A(n13235), .B(n13272), .C(n13350), .D(n10809), .Y(n13869)
         );
  INVX1 U9447 ( .A(n12338), .Y(n12365) );
  AOI22X1 U9448 ( .A(\lamb/scale_ds1/genblk1[1].mult/added[1] ), .B(n11053), 
        .C(n12365), .D(n10754), .Y(n12342) );
  AOI21X1 U9449 ( .A(n12342), .B(n12341), .C(n10465), .Y(n12348) );
  OAI21X1 U9450 ( .A(n12345), .B(n12343), .C(n12344), .Y(n12346) );
  NAND2X1 U9451 ( .A(n11147), .B(n12346), .Y(n12347) );
  HAX1 U9452 ( .A(n12348), .B(n12347), .YS(n13935) );
  AOI22X1 U9453 ( .A(n11227), .B(n10732), .C(n13935), .D(n13841), .Y(n13039)
         );
  INVX1 U9454 ( .A(n10471), .Y(n13274) );
  AOI22X1 U9455 ( .A(n13235), .B(n13274), .C(n13348), .D(n10809), .Y(n13178)
         );
  AOI21X1 U9456 ( .A(n10653), .B(n12350), .C(n12349), .Y(n12352) );
  AOI22X1 U9457 ( .A(\lamb/scale_ts1/genblk1[1].mult/added[1] ), .B(n12355), 
        .C(\lamb/scale_ts1/genblk1[1].mult/added[2] ), .D(n12354), .Y(n12359)
         );
  INVX1 U9458 ( .A(n11147), .Y(n12357) );
  AOI21X1 U9459 ( .A(n12359), .B(n11057), .C(n12357), .Y(n12370) );
  INVX1 U9460 ( .A(n10631), .Y(n12362) );
  AOI22X1 U9461 ( .A(\lamb/scale_ds1/genblk1[1].mult/added[1] ), .B(n12365), 
        .C(n12364), .D(n10950), .Y(n12368) );
  AOI21X1 U9462 ( .A(n12368), .B(n12367), .C(n10465), .Y(n12369) );
  HAX1 U9463 ( .A(n12370), .B(n12369), .YS(n13934) );
  INVX1 U9464 ( .A(n13934), .Y(n13200) );
  AOI22X1 U9465 ( .A(n11227), .B(n10817), .C(n13200), .D(n13841), .Y(n13045)
         );
  AOI21X1 U9466 ( .A(n10733), .B(n10658), .C(n10690), .Y(n13036) );
  INVX1 U9467 ( .A(n10676), .Y(n12371) );
  AOI21X1 U9468 ( .A(n13037), .B(n10431), .C(n12371), .Y(n12396) );
  OAI21X1 U9469 ( .A(n12376), .B(n12372), .C(n11099), .Y(n12373) );
  HAX1 U9470 ( .A(n12374), .B(n12373), .YS(n13011) );
  NOR3X1 U9471 ( .A(n12289), .B(n10634), .C(
        \lamb/scale_ts3/genblk1[2].mult/added[3] ), .Y(n12411) );
  INVX1 U9472 ( .A(n12376), .Y(n12377) );
  OAI21X1 U9473 ( .A(\lamb/scale_ts3/genblk1[2].mult/added[1] ), .B(n12411), 
        .C(n12377), .Y(n12378) );
  INVX1 U9474 ( .A(n11099), .Y(n12412) );
  AOI21X1 U9475 ( .A(n12379), .B(n12378), .C(n12412), .Y(n12385) );
  NOR3X1 U9476 ( .A(\lamb/scale_ds3/genblk1[2].mult/added[3] ), .B(n12380), 
        .C(n12178), .Y(n12418) );
  OAI21X1 U9477 ( .A(n12418), .B(\lamb/scale_ds3/genblk1[2].mult/added[1] ), 
        .C(n11018), .Y(n12382) );
  NAND2X1 U9478 ( .A(n12383), .B(n12382), .Y(n12416) );
  NAND2X1 U9479 ( .A(n12416), .B(n11155), .Y(n12384) );
  HAX1 U9480 ( .A(n12385), .B(n12384), .YS(n12633) );
  OAI21X1 U9481 ( .A(n11182), .B(n12386), .C(n10516), .Y(n12388) );
  AOI22X1 U9482 ( .A(\lamb/scale_ts3/genblk1[2].mult/added[2] ), .B(n12411), 
        .C(n10428), .D(n12388), .Y(n12393) );
  INVX1 U9483 ( .A(\lamb/scale_ts3/genblk1[2].mult/added[2] ), .Y(n12390) );
  NAND3X1 U9484 ( .A(\lamb/scale_ts3/genblk1[2].mult/added[1] ), .B(n12392), 
        .C(n11087), .Y(n12413) );
  NAND3X1 U9485 ( .A(n12394), .B(n12393), .C(n10408), .Y(n12395) );
  NAND2X1 U9486 ( .A(n11099), .B(n12395), .Y(n12406) );
  AOI22X1 U9487 ( .A(\lamb/scale_ds3/genblk1[2].mult/added[2] ), .B(n12418), 
        .C(n12417), .D(n12397), .Y(n12403) );
  INVX1 U9488 ( .A(n12398), .Y(n12399) );
  OAI21X1 U9489 ( .A(n12400), .B(\lamb/scale_ds3/genblk1[2].mult/added[2] ), 
        .C(n12399), .Y(n12401) );
  NAND3X1 U9490 ( .A(n10923), .B(n10433), .C(n10436), .Y(n12404) );
  XNOR2X1 U9491 ( .A(n12406), .B(n10390), .Y(n13015) );
  NAND2X1 U9492 ( .A(n11019), .B(n13015), .Y(n12634) );
  INVX1 U9493 ( .A(n13011), .Y(n12627) );
  NAND2X1 U9494 ( .A(n12408), .B(n10516), .Y(n12409) );
  AOI22X1 U9495 ( .A(\lamb/scale_ts3/genblk1[2].mult/added[1] ), .B(n12411), 
        .C(n11087), .D(n12409), .Y(n12414) );
  AOI21X1 U9496 ( .A(n12414), .B(n10408), .C(n12412), .Y(n12426) );
  INVX1 U9497 ( .A(n12415), .Y(n12424) );
  INVX1 U9498 ( .A(n12416), .Y(n12421) );
  AOI22X1 U9499 ( .A(\lamb/scale_ds3/genblk1[2].mult/added[1] ), .B(n12418), 
        .C(\lamb/scale_ds3/genblk1[2].mult/added[2] ), .D(n12417), .Y(n12419)
         );
  OAI21X1 U9500 ( .A(n12421), .B(n10436), .C(n12419), .Y(n12423) );
  OAI21X1 U9501 ( .A(n12424), .B(n12423), .C(n11155), .Y(n12425) );
  HAX1 U9502 ( .A(n12426), .B(n12425), .YS(n13013) );
  OAI21X1 U9503 ( .A(n10750), .B(n12633), .C(n13013), .Y(n13009) );
  NOR2X1 U9504 ( .A(n12634), .B(n13009), .Y(n12842) );
  AOI21X1 U9505 ( .A(n13002), .B(n12994), .C(n12842), .Y(n12602) );
  INVX1 U9506 ( .A(\forney/pe0/mult0/added [1]), .Y(n12570) );
  OR2X1 U9507 ( .A(\forney/pe0/mult0/added [4]), .B(\add_x_87/n1 ), .Y(n12535)
         );
  INVX1 U9508 ( .A(n12535), .Y(n12427) );
  INVX1 U9509 ( .A(\forney/pe0/mult0/added [3]), .Y(n12530) );
  AOI22X1 U9510 ( .A(\forney/pe0/mult0/added [3]), .B(n12427), .C(n12572), .D(
        n12530), .Y(n12532) );
  OAI21X1 U9511 ( .A(n12570), .B(n12532), .C(n10661), .Y(n12428) );
  INVX1 U9512 ( .A(\forney/pe0/mult0/added [2]), .Y(n12536) );
  NAND2X1 U9513 ( .A(\forney/pe0/mult0/added [2]), .B(
        \forney/pe0/mult0/added [1]), .Y(n12533) );
  INVX1 U9514 ( .A(n12533), .Y(n12429) );
  NOR3X1 U9515 ( .A(\forney/pe0/mult0/added [3]), .B(
        \forney/pe0/mult0/added [4]), .C(\add_x_87/n1 ), .Y(n12569) );
  AOI21X1 U9516 ( .A(n12429), .B(n10661), .C(n12569), .Y(n12575) );
  NAND3X1 U9517 ( .A(\forney/pe0/mult0/added [3]), .B(n12535), .C(n12570), .Y(
        n12600) );
  OR2X1 U9518 ( .A(n12536), .B(n12600), .Y(n12571) );
  NAND3X1 U9519 ( .A(n11059), .B(n10405), .C(n12571), .Y(n12430) );
  NAND2X1 U9520 ( .A(n11148), .B(n12430), .Y(n12529) );
  NAND2X1 U9521 ( .A(n13903), .B(n13893), .Y(n12863) );
  INVX1 U9522 ( .A(n12863), .Y(n13693) );
  NAND2X1 U9523 ( .A(n13888), .B(n12431), .Y(n12789) );
  OR2X1 U9524 ( .A(n12833), .B(n12789), .Y(n12857) );
  OR2X1 U9525 ( .A(n12856), .B(n12857), .Y(n12432) );
  INVX1 U9526 ( .A(n12862), .Y(n13387) );
  NAND3X1 U9527 ( .A(\lamb/scale_ds3/genblk1[3].mult/added[3] ), .B(
        \add_x_120/n1 ), .C(\lamb/scale_ds3/genblk1[3].mult/added[4] ), .Y(
        n12434) );
  INVX1 U9528 ( .A(n12434), .Y(n12584) );
  NAND2X1 U9529 ( .A(n12584), .B(n11193), .Y(n12544) );
  INVX1 U9530 ( .A(\lamb/scale_ds3/genblk1[3].mult/added[1] ), .Y(n12546) );
  AOI21X1 U9531 ( .A(\add_x_120/n1 ), .B(
        \lamb/scale_ds3/genblk1[3].mult/added[4] ), .C(
        \lamb/scale_ds3/genblk1[3].mult/added[3] ), .Y(n12543) );
  INVX1 U9532 ( .A(n10537), .Y(n12433) );
  OR2X1 U9533 ( .A(\add_x_120/n1 ), .B(
        \lamb/scale_ds3/genblk1[3].mult/added[4] ), .Y(n12547) );
  NOR2X1 U9534 ( .A(n12546), .B(n11130), .Y(n12611) );
  INVX1 U9535 ( .A(n12611), .Y(n12435) );
  NOR3X1 U9536 ( .A(\lamb/scale_ds3/genblk1[3].mult/added[3] ), .B(
        \add_x_120/n1 ), .C(\lamb/scale_ds3/genblk1[3].mult/added[4] ), .Y(
        n12437) );
  OAI21X1 U9537 ( .A(n12549), .B(n12437), .C(n12434), .Y(n12585) );
  NAND3X1 U9538 ( .A(n12544), .B(n12435), .C(n12585), .Y(n12510) );
  AND2X1 U9539 ( .A(\add_x_120/n1 ), .B(
        \lamb/scale_ds3/genblk1[3].mult/added[4] ), .Y(n12436) );
  NOR3X1 U9540 ( .A(\lamb/scale_ds3/genblk1[3].mult/added[1] ), .B(n12436), 
        .C(n10667), .Y(n12612) );
  OAI21X1 U9541 ( .A(n12612), .B(n12437), .C(
        \lamb/scale_ds3/genblk1[3].mult/added[2] ), .Y(n12586) );
  INVX1 U9542 ( .A(n12586), .Y(n12509) );
  INVX1 U9543 ( .A(n10444), .Y(n13868) );
  INVX1 U9544 ( .A(n10726), .Y(n12690) );
  INVX1 U9545 ( .A(n10732), .Y(n12691) );
  AOI21X1 U9546 ( .A(n12691), .B(n10549), .C(n10816), .Y(n13172) );
  AOI21X1 U9547 ( .A(n10425), .B(n10432), .C(n12438), .Y(n12495) );
  INVX1 U9548 ( .A(\lamb/scale_ts2/genblk1[2].mult/added[3] ), .Y(n12439) );
  NOR2X1 U9549 ( .A(\add_x_130/n1 ), .B(
        \lamb/scale_ts2/genblk1[2].mult/added[4] ), .Y(n12460) );
  NAND2X1 U9550 ( .A(\add_x_130/n1 ), .B(
        \lamb/scale_ts2/genblk1[2].mult/added[4] ), .Y(n12445) );
  NAND2X1 U9551 ( .A(n12439), .B(n12445), .Y(n12440) );
  INVX1 U9552 ( .A(\lamb/scale_ts2/genblk1[2].mult/added[1] ), .Y(n12441) );
  NAND3X1 U9553 ( .A(\add_x_130/n1 ), .B(
        \lamb/scale_ts2/genblk1[2].mult/added[4] ), .C(
        \lamb/scale_ts2/genblk1[2].mult/added[3] ), .Y(n12444) );
  OAI21X1 U9554 ( .A(n10993), .B(n12441), .C(n12444), .Y(n12443) );
  NOR2X1 U9555 ( .A(\lamb/scale_ts2/genblk1[2].mult/added[1] ), .B(n12462), 
        .Y(n12446) );
  NAND2X1 U9556 ( .A(\lamb/scale_ts2/genblk1[2].mult/added[2] ), .B(n11013), 
        .Y(n12442) );
  OAI21X1 U9557 ( .A(\lamb/scale_ts2/genblk1[2].mult/added[2] ), .B(n12443), 
        .C(n12442), .Y(n12487) );
  NOR3X1 U9558 ( .A(\add_x_130/n1 ), .B(
        \lamb/scale_ts2/genblk1[2].mult/added[4] ), .C(
        \lamb/scale_ts2/genblk1[2].mult/added[3] ), .Y(n12485) );
  OAI21X1 U9559 ( .A(n12485), .B(n12483), .C(n12444), .Y(n12484) );
  INVX1 U9560 ( .A(n12445), .Y(n12459) );
  NAND3X1 U9561 ( .A(n12446), .B(n12459), .C(
        \lamb/scale_ts2/genblk1[2].mult/added[2] ), .Y(n12464) );
  NAND3X1 U9562 ( .A(n12487), .B(n12484), .C(n10434), .Y(n12447) );
  NAND2X1 U9563 ( .A(n11149), .B(n12447), .Y(n12458) );
  OR2X1 U9564 ( .A(\add_x_134/n1 ), .B(
        \lamb/scale_ds2/genblk1[2].mult/added[4] ), .Y(n12448) );
  NAND2X1 U9565 ( .A(\add_x_134/n1 ), .B(
        \lamb/scale_ds2/genblk1[2].mult/added[4] ), .Y(n12451) );
  INVX1 U9566 ( .A(n12451), .Y(n12468) );
  NAND2X1 U9567 ( .A(\lamb/scale_ds2/genblk1[2].mult/added[3] ), .B(n12448), 
        .Y(n12469) );
  NOR2X1 U9568 ( .A(\lamb/scale_ds2/genblk1[2].mult/added[1] ), .B(n12469), 
        .Y(n12452) );
  NAND2X1 U9569 ( .A(\lamb/scale_ds2/genblk1[2].mult/added[2] ), .B(n12481), 
        .Y(n12471) );
  NAND3X1 U9570 ( .A(n12468), .B(n12452), .C(n11090), .Y(n12472) );
  NAND3X1 U9571 ( .A(\add_x_134/n1 ), .B(
        \lamb/scale_ds2/genblk1[2].mult/added[4] ), .C(
        \lamb/scale_ds2/genblk1[2].mult/added[3] ), .Y(n12450) );
  NAND3X1 U9572 ( .A(\lamb/scale_ds2/genblk1[2].mult/added[2] ), .B(
        \lamb/scale_ds2/genblk1[2].mult/added[1] ), .C(n12450), .Y(n12478) );
  NAND3X1 U9573 ( .A(n12481), .B(n10406), .C(n12478), .Y(n12456) );
  INVX1 U9574 ( .A(\lamb/scale_ds2/genblk1[2].mult/added[3] ), .Y(n12449) );
  INVX1 U9575 ( .A(n12448), .Y(n12467) );
  AOI22X1 U9576 ( .A(n12468), .B(n12449), .C(n12467), .D(
        \lamb/scale_ds2/genblk1[2].mult/added[3] ), .Y(n12499) );
  INVX1 U9577 ( .A(n12450), .Y(n12454) );
  NAND2X1 U9578 ( .A(n12452), .B(n12451), .Y(n12504) );
  OAI21X1 U9579 ( .A(\lamb/scale_ds2/genblk1[2].mult/added[2] ), .B(n12454), 
        .C(n12453), .Y(n12480) );
  OAI21X1 U9580 ( .A(n10558), .B(n11091), .C(n12480), .Y(n12455) );
  NOR2X1 U9581 ( .A(n13933), .B(n13937), .Y(n13201) );
  INVX1 U9582 ( .A(n13935), .Y(n13205) );
  NAND2X1 U9583 ( .A(n13933), .B(n13937), .Y(n13199) );
  AOI21X1 U9584 ( .A(n13205), .B(n13199), .C(n13934), .Y(n13202) );
  OAI21X1 U9585 ( .A(n12456), .B(n12455), .C(n11154), .Y(n12457) );
  HAX1 U9586 ( .A(n12458), .B(n12457), .YS(n13053) );
  NOR3X1 U9587 ( .A(n12460), .B(\lamb/scale_ts2/genblk1[2].mult/added[3] ), 
        .C(n12459), .Y(n12491) );
  AOI22X1 U9588 ( .A(\lamb/scale_ts2/genblk1[2].mult/added[2] ), .B(n12491), 
        .C(n12461), .D(n10645), .Y(n12465) );
  OR2X1 U9589 ( .A(\lamb/scale_ts2/genblk1[2].mult/added[2] ), .B(n12462), .Y(
        n12493) );
  OAI21X1 U9590 ( .A(n12485), .B(n10930), .C(
        \lamb/scale_ts2/genblk1[2].mult/added[1] ), .Y(n12463) );
  NAND3X1 U9591 ( .A(n12465), .B(n10434), .C(n12463), .Y(n12466) );
  NAND2X1 U9592 ( .A(n11149), .B(n12466), .Y(n12477) );
  AOI21X1 U9593 ( .A(\lamb/scale_ds2/genblk1[2].mult/added[2] ), .B(
        \lamb/scale_ds2/genblk1[2].mult/added[1] ), .C(n10558), .Y(n12475) );
  NOR3X1 U9594 ( .A(n12468), .B(n12467), .C(
        \lamb/scale_ds2/genblk1[2].mult/added[3] ), .Y(n12501) );
  AOI22X1 U9595 ( .A(\lamb/scale_ds2/genblk1[2].mult/added[1] ), .B(n10628), 
        .C(\lamb/scale_ds2/genblk1[2].mult/added[2] ), .D(n12501), .Y(n12473)
         );
  NAND2X1 U9596 ( .A(n10877), .B(n12469), .Y(n12470) );
  NAND3X1 U9597 ( .A(n12473), .B(n10406), .C(n12502), .Y(n12474) );
  OAI21X1 U9598 ( .A(n12475), .B(n12474), .C(n11154), .Y(n12476) );
  HAX1 U9599 ( .A(n12477), .B(n12476), .YS(n13061) );
  NOR2X1 U9600 ( .A(n13053), .B(n13061), .Y(n13058) );
  OAI21X1 U9601 ( .A(\lamb/scale_ds2/genblk1[2].mult/added[1] ), .B(n12501), 
        .C(n12478), .Y(n12479) );
  AOI22X1 U9602 ( .A(n10628), .B(n10877), .C(n12480), .D(n12479), .Y(n12482)
         );
  NAND2X1 U9603 ( .A(n12482), .B(n11154), .Y(n12490) );
  AOI22X1 U9604 ( .A(\lamb/scale_ts2/genblk1[2].mult/added[1] ), .B(n12484), 
        .C(n12491), .D(n10645), .Y(n12486) );
  NAND2X1 U9605 ( .A(\lamb/scale_ts2/genblk1[2].mult/added[2] ), .B(n12485), 
        .Y(n12492) );
  NAND3X1 U9606 ( .A(n12487), .B(n12486), .C(n12492), .Y(n12488) );
  NAND2X1 U9607 ( .A(n11149), .B(n12488), .Y(n12489) );
  HAX1 U9608 ( .A(n12490), .B(n12489), .YS(n12719) );
  AOI22X1 U9609 ( .A(\lamb/scale_ts2/genblk1[2].mult/added[1] ), .B(n12494), 
        .C(\lamb/scale_ts2/genblk1[2].mult/added[2] ), .D(n12461), .Y(n12497)
         );
  INVX1 U9610 ( .A(n11149), .Y(n12496) );
  AOI21X1 U9611 ( .A(n11013), .B(n12497), .C(n12496), .Y(n12508) );
  INVX1 U9612 ( .A(n10558), .Y(n12500) );
  AOI22X1 U9613 ( .A(\lamb/scale_ds2/genblk1[2].mult/added[1] ), .B(n12501), 
        .C(\lamb/scale_ds2/genblk1[2].mult/added[2] ), .D(n12500), .Y(n12503)
         );
  NAND3X1 U9614 ( .A(n12504), .B(n12503), .C(n12502), .Y(n12506) );
  NAND2X1 U9615 ( .A(n12506), .B(n11154), .Y(n12507) );
  HAX1 U9616 ( .A(n12508), .B(n12507), .YS(n13064) );
  INVX1 U9617 ( .A(n13064), .Y(n12720) );
  AOI21X1 U9618 ( .A(n12719), .B(n10651), .C(n12720), .Y(n13057) );
  OAI21X1 U9619 ( .A(n12510), .B(n12509), .C(n11146), .Y(n12527) );
  INVX1 U9620 ( .A(n13876), .Y(n13191) );
  AOI22X1 U9621 ( .A(n11227), .B(n12511), .C(n13191), .D(n13841), .Y(n12624)
         );
  AOI22X1 U9622 ( .A(n11227), .B(n13154), .C(n13880), .D(n13841), .Y(n13025)
         );
  INVX1 U9623 ( .A(n13157), .Y(n13152) );
  AOI22X1 U9624 ( .A(n11227), .B(n13152), .C(n13879), .D(n13841), .Y(n13028)
         );
  INVX1 U9625 ( .A(n10678), .Y(n12512) );
  INVX1 U9626 ( .A(n13194), .Y(n13193) );
  AOI22X1 U9627 ( .A(n11227), .B(n13158), .C(n13193), .D(n13841), .Y(n12513)
         );
  AOI22X1 U9628 ( .A(n10543), .B(n10813), .C(n12512), .D(n12513), .Y(n12626)
         );
  INVX1 U9629 ( .A(n12513), .Y(n13027) );
  NOR2X1 U9630 ( .A(n10543), .B(n13034), .Y(n13023) );
  OAI21X1 U9631 ( .A(n13027), .B(n10812), .C(n13023), .Y(n13031) );
  OAI21X1 U9632 ( .A(n12626), .B(n13031), .C(n10676), .Y(n12607) );
  INVX1 U9633 ( .A(n12607), .Y(n12564) );
  NAND3X1 U9634 ( .A(\add_x_116/n1 ), .B(
        \lamb/scale_ts3/genblk1[3].mult/added[4] ), .C(
        \lamb/scale_ts3/genblk1[3].mult/added[3] ), .Y(n12520) );
  INVX1 U9635 ( .A(n10561), .Y(n12515) );
  INVX1 U9636 ( .A(\lamb/scale_ts3/genblk1[3].mult/added[1] ), .Y(n12518) );
  NAND3X1 U9637 ( .A(\lamb/scale_ts3/genblk1[3].mult/added[2] ), .B(n12515), 
        .C(n12518), .Y(n12560) );
  INVX1 U9638 ( .A(n10522), .Y(n12552) );
  NOR3X1 U9639 ( .A(\add_x_116/n1 ), .B(
        \lamb/scale_ts3/genblk1[3].mult/added[4] ), .C(
        \lamb/scale_ts3/genblk1[3].mult/added[3] ), .Y(n12554) );
  AOI21X1 U9640 ( .A(n12552), .B(n10561), .C(n12554), .Y(n12580) );
  NOR2X1 U9641 ( .A(\add_x_116/n1 ), .B(
        \lamb/scale_ts3/genblk1[3].mult/added[4] ), .Y(n12519) );
  INVX1 U9642 ( .A(n12519), .Y(n12517) );
  NAND2X1 U9643 ( .A(\add_x_116/n1 ), .B(
        \lamb/scale_ts3/genblk1[3].mult/added[4] ), .Y(n12516) );
  INVX1 U9644 ( .A(\lamb/scale_ts3/genblk1[3].mult/added[3] ), .Y(n12558) );
  AOI22X1 U9645 ( .A(\lamb/scale_ts3/genblk1[3].mult/added[3] ), .B(n12517), 
        .C(n12516), .D(n12558), .Y(n12605) );
  NAND2X1 U9646 ( .A(n10522), .B(n12605), .Y(n12562) );
  INVX1 U9647 ( .A(n12562), .Y(n12524) );
  NAND2X1 U9648 ( .A(\lamb/scale_ts3/genblk1[3].mult/added[2] ), .B(n12518), 
        .Y(n12522) );
  AOI21X1 U9649 ( .A(\lamb/scale_ts3/genblk1[3].mult/added[4] ), .B(
        \add_x_116/n1 ), .C(n12519), .Y(n12557) );
  NAND2X1 U9650 ( .A(\lamb/scale_ts3/genblk1[3].mult/added[3] ), .B(n12557), 
        .Y(n12553) );
  OR2X1 U9651 ( .A(\lamb/scale_ts3/genblk1[3].mult/added[2] ), .B(n10561), .Y(
        n12556) );
  INVX1 U9652 ( .A(n12556), .Y(n12521) );
  AOI21X1 U9653 ( .A(\lamb/scale_ts3/genblk1[3].mult/added[2] ), .B(n12554), 
        .C(n12521), .Y(n12604) );
  OAI21X1 U9654 ( .A(n12522), .B(n12553), .C(n12604), .Y(n12523) );
  AOI21X1 U9655 ( .A(\lamb/scale_ts3/genblk1[3].mult/added[1] ), .B(n12524), 
        .C(n12523), .Y(n12582) );
  NAND3X1 U9656 ( .A(n12560), .B(n10394), .C(n11081), .Y(n12525) );
  NAND2X1 U9657 ( .A(n12564), .B(n12525), .Y(n12526) );
  HAX1 U9658 ( .A(n12527), .B(n12526), .YS(n12873) );
  XNOR2X1 U9659 ( .A(n12529), .B(n10391), .Y(n12951) );
  NAND3X1 U9660 ( .A(n12530), .B(n12535), .C(n11132), .Y(n12595) );
  OAI21X1 U9661 ( .A(\forney/pe0/mult0/added [1]), .B(n10661), .C(n10597), .Y(
        n12534) );
  INVX1 U9662 ( .A(n12532), .Y(n12598) );
  AOI22X1 U9663 ( .A(\forney/pe0/mult0/added [2]), .B(n12534), .C(n12598), .D(
        n12533), .Y(n12540) );
  NAND3X1 U9664 ( .A(\forney/pe0/mult0/added [3]), .B(n12536), .C(n12535), .Y(
        n12594) );
  INVX1 U9665 ( .A(n12594), .Y(n12537) );
  OAI21X1 U9666 ( .A(n12569), .B(n12537), .C(\forney/pe0/mult0/added [1]), .Y(
        n12539) );
  INVX1 U9667 ( .A(n11148), .Y(n12538) );
  AOI21X1 U9668 ( .A(n10925), .B(n12539), .C(n12538), .Y(n12568) );
  INVX1 U9669 ( .A(\lamb/scale_ds3/genblk1[3].mult/added[2] ), .Y(n12583) );
  AOI22X1 U9670 ( .A(n12583), .B(n10667), .C(n12546), .D(n11130), .Y(n12542)
         );
  OAI21X1 U9671 ( .A(n10537), .B(n11193), .C(n12542), .Y(n12615) );
  AND2X1 U9672 ( .A(n10537), .B(n12547), .Y(n12610) );
  NAND2X1 U9673 ( .A(n12610), .B(n11193), .Y(n12588) );
  NAND2X1 U9674 ( .A(n12544), .B(n12588), .Y(n12550) );
  OAI21X1 U9675 ( .A(n12547), .B(n12546), .C(n11130), .Y(n12548) );
  AOI22X1 U9676 ( .A(\lamb/scale_ds3/genblk1[3].mult/added[2] ), .B(n12550), 
        .C(n11193), .D(n12548), .Y(n12551) );
  AOI21X1 U9677 ( .A(n12615), .B(n12551), .C(n12616), .Y(n12566) );
  OR2X1 U9678 ( .A(n12553), .B(n12552), .Y(n12608) );
  INVX1 U9679 ( .A(n12554), .Y(n12555) );
  NAND3X1 U9680 ( .A(n12608), .B(n12556), .C(n12555), .Y(n12559) );
  AOI22X1 U9681 ( .A(\lamb/scale_ts3/genblk1[3].mult/added[1] ), .B(n12559), 
        .C(\lamb/scale_ts3/genblk1[3].mult/added[2] ), .D(n12603), .Y(n12561)
         );
  NAND3X1 U9682 ( .A(n12562), .B(n12561), .C(n12560), .Y(n12563) );
  XNOR2X1 U9683 ( .A(n12566), .B(n10983), .Y(n12904) );
  NAND2X1 U9684 ( .A(n11157), .B(n12904), .Y(n12567) );
  HAX1 U9685 ( .A(n12568), .B(n12567), .YS(n12954) );
  NAND2X1 U9686 ( .A(n12951), .B(n12954), .Y(n13479) );
  NAND2X1 U9687 ( .A(\forney/pe0/mult0/added [2]), .B(n12569), .Y(n12596) );
  NAND2X1 U9688 ( .A(n12570), .B(n10597), .Y(n12574) );
  INVX1 U9689 ( .A(n12571), .Y(n12573) );
  AOI22X1 U9690 ( .A(n10405), .B(n12574), .C(n12573), .D(n11132), .Y(n12577)
         );
  NAND3X1 U9691 ( .A(n12596), .B(n12577), .C(n11059), .Y(n12578) );
  NAND2X1 U9692 ( .A(n11148), .B(n12578), .Y(n12593) );
  AOI22X1 U9693 ( .A(\lamb/scale_ts3/genblk1[3].mult/added[1] ), .B(n10394), 
        .C(n12603), .D(n10522), .Y(n12581) );
  AOI21X1 U9694 ( .A(n11081), .B(n12581), .C(n12607), .Y(n12591) );
  AOI22X1 U9695 ( .A(\lamb/scale_ds3/genblk1[3].mult/added[1] ), .B(n12585), 
        .C(n12584), .D(n12583), .Y(n12587) );
  NAND3X1 U9696 ( .A(n12588), .B(n12587), .C(n12586), .Y(n12589) );
  XNOR2X1 U9697 ( .A(n12591), .B(n10392), .Y(n12867) );
  NAND2X1 U9698 ( .A(n12867), .B(n11157), .Y(n12592) );
  HAX1 U9699 ( .A(n12593), .B(n12592), .YS(n12952) );
  NAND3X1 U9700 ( .A(n12596), .B(n10597), .C(n12594), .Y(n12597) );
  AOI22X1 U9701 ( .A(\forney/pe0/mult0/added [2]), .B(n12598), .C(
        \forney/pe0/mult0/added [1]), .D(n12597), .Y(n12599) );
  OAI21X1 U9702 ( .A(n12600), .B(n12572), .C(n12599), .Y(n12601) );
  NAND2X1 U9703 ( .A(n11148), .B(n12601), .Y(n12622) );
  NAND2X1 U9704 ( .A(n12604), .B(n10985), .Y(n12606) );
  AOI22X1 U9705 ( .A(\lamb/scale_ts3/genblk1[3].mult/added[1] ), .B(n12606), 
        .C(\lamb/scale_ts3/genblk1[3].mult/added[2] ), .D(n12605), .Y(n12609)
         );
  AOI21X1 U9706 ( .A(n12609), .B(n12608), .C(n12607), .Y(n12619) );
  AOI22X1 U9707 ( .A(\lamb/scale_ds3/genblk1[3].mult/added[2] ), .B(n12611), 
        .C(\lamb/scale_ds3/genblk1[3].mult/added[1] ), .D(n12610), .Y(n12614)
         );
  INVX1 U9708 ( .A(n12612), .Y(n12613) );
  NAND3X1 U9709 ( .A(n12615), .B(n12614), .C(n12613), .Y(n12617) );
  XNOR2X1 U9710 ( .A(n10982), .B(n10393), .Y(n12887) );
  NAND2X1 U9711 ( .A(n12887), .B(n11157), .Y(n12621) );
  HAX1 U9712 ( .A(n12622), .B(n12621), .YS(n12717) );
  INVX1 U9713 ( .A(n12717), .Y(n12955) );
  NAND2X1 U9714 ( .A(n12952), .B(n12955), .Y(n12714) );
  OR2X1 U9715 ( .A(n12951), .B(n12954), .Y(n12953) );
  INVX1 U9716 ( .A(n12953), .Y(n12715) );
  NAND2X1 U9717 ( .A(n12717), .B(n11165), .Y(n12713) );
  OAI21X1 U9718 ( .A(n12714), .B(n12715), .C(n12713), .Y(n12623) );
  AND2X1 U9719 ( .A(n13479), .B(n12623), .Y(\forney/m0/logB [1]) );
  NAND2X1 U9720 ( .A(n10678), .B(n13027), .Y(n13022) );
  INVX1 U9721 ( .A(n13022), .Y(n13024) );
  OAI21X1 U9722 ( .A(n10743), .B(n13024), .C(n10812), .Y(n12625) );
  AND2X1 U9723 ( .A(n12626), .B(n12625), .Y(
        \lamb/scale_ts3/genblk1[3].mult/logA[1] ) );
  INVX1 U9724 ( .A(n12633), .Y(n13008) );
  NAND2X1 U9725 ( .A(n12627), .B(n13008), .Y(n12635) );
  AOI21X1 U9726 ( .A(n11019), .B(n12635), .C(n13013), .Y(n12629) );
  AOI21X1 U9727 ( .A(n12630), .B(n10659), .C(n10576), .Y(n12632) );
  INVX1 U9728 ( .A(n12631), .Y(n13004) );
  OR2X1 U9729 ( .A(n12632), .B(n13004), .Y(\forney/pe0/mult0/logB [0]) );
  NAND2X1 U9730 ( .A(n10750), .B(n12633), .Y(n13018) );
  AOI21X1 U9731 ( .A(n12634), .B(n13018), .C(n13013), .Y(n12636) );
  INVX1 U9732 ( .A(n12635), .Y(n13014) );
  OR2X1 U9733 ( .A(n12636), .B(n13014), .Y(\forney/pe0/mult0/logA [3]) );
  MUX2X1 U9734 ( .B(n12639), .A(n12638), .S(n12637), .Y(n12655) );
  MUX2X1 U9735 ( .B(n11145), .A(n12641), .S(n12640), .Y(n12643) );
  MUX2X1 U9736 ( .B(n12645), .A(n12644), .S(n12643), .Y(n12654) );
  AOI22X1 U9737 ( .A(msg[28]), .B(msg[48]), .C(n12646), .D(n13717), .Y(n12648)
         );
  AOI22X1 U9738 ( .A(msg[8]), .B(msg[13]), .C(n13764), .D(n13787), .Y(n12647)
         );
  FAX1 U9739 ( .A(n12649), .B(n10755), .C(n10696), .YS(n12650) );
  MUX2X1 U9740 ( .B(n11167), .A(n12651), .S(n12650), .Y(n12653) );
  FAX1 U9741 ( .A(n12655), .B(n12654), .C(n12653), .YS(n12656) );
  MUX2X1 U9742 ( .B(n12658), .A(n12657), .S(n12656), .Y(n12661) );
  OAI21X1 U9743 ( .A(n12670), .B(n12661), .C(n11133), .Y(
        \lamb/scale_ts0/genblk1[0].mult/logA[0] ) );
  AND2X1 U9744 ( .A(n10851), .B(\lamb/scale_ts0/genblk1[0].mult/logA[0] ), .Y(
        \lamb/scale_ts1/genblk1[0].mult/logA[0] ) );
  AOI21X1 U9745 ( .A(n12664), .B(n12665), .C(n12659), .Y(n12662) );
  AOI22X1 U9746 ( .A(n12667), .B(n12662), .C(n12661), .D(n10957), .Y(
        \lamb/scale_ts0/genblk1[0].mult/logA[3] ) );
  AOI21X1 U9747 ( .A(n12665), .B(n12664), .C(n12663), .Y(n12666) );
  MUX2X1 U9748 ( .B(n11133), .A(n12667), .S(n12666), .Y(n12669) );
  AOI21X1 U9749 ( .A(n12671), .B(n12670), .C(n12669), .Y(
        \lamb/scale_ts0/genblk1[0].mult/logA[2] ) );
  AND2X1 U9750 ( .A(n10851), .B(n10786), .Y(
        \lamb/scale_ts1/genblk1[0].mult/logA[2] ) );
  AND2X1 U9751 ( .A(n10851), .B(n10787), .Y(
        \lamb/scale_ts1/genblk1[0].mult/logA[1] ) );
  AND2X1 U9752 ( .A(\lamb/scale_ts1/genblk1[3].mult/logA[0] ), .B(n13841), .Y(
        \lamb/scale_bs3/genblk1[0].mult/logA[0] ) );
  OAI21X1 U9753 ( .A(n12675), .B(n11010), .C(n12674), .Y(n12676) );
  AOI21X1 U9754 ( .A(n11010), .B(n12677), .C(n12676), .Y(n10377) );
  AND2X1 U9755 ( .A(n10701), .B(n12682), .Y(
        \lamb/scale_ls2/genblk1[1].mult/logA[3] ) );
  AND2X1 U9756 ( .A(\lamb/scale_ls2/genblk1[1].mult/logA[3] ), .B(n13841), .Y(
        \lamb/scale_bs3/genblk1[0].mult/logA[3] ) );
  AND2X1 U9757 ( .A(\lamb/scale_ls2/genblk1[1].mult/logA[2] ), .B(n13841), .Y(
        \lamb/scale_bs3/genblk1[0].mult/logA[2] ) );
  NAND2X1 U9758 ( .A(n12679), .B(n10689), .Y(n12681) );
  AOI21X1 U9759 ( .A(n12681), .B(n11124), .C(n12680), .Y(n10378) );
  AND2X1 U9760 ( .A(n10792), .B(n12682), .Y(n10372) );
  AND2X1 U9761 ( .A(n10372), .B(n13841), .Y(
        \lamb/scale_bs3/genblk1[0].mult/logA[1] ) );
  AND2X1 U9762 ( .A(n13258), .B(n10379), .Y(
        \lamb/scale_ls2/genblk1[0].mult/logA[0] ) );
  AND2X1 U9763 ( .A(n10851), .B(n10701), .Y(
        \lamb/scale_ls2/genblk1[0].mult/logA[3] ) );
  AND2X1 U9764 ( .A(n10851), .B(n10792), .Y(
        \lamb/scale_ls2/genblk1[0].mult/logA[1] ) );
  INVX1 U9765 ( .A(n10528), .Y(n12688) );
  OAI21X1 U9766 ( .A(n13083), .B(n10749), .C(n13845), .Y(n10376) );
  AND2X1 U9767 ( .A(n13224), .B(n10376), .Y(
        \lamb/scale_bs2/genblk1[0].mult/logA[0] ) );
  NAND3X1 U9768 ( .A(n13229), .B(n10818), .C(n10749), .Y(n12687) );
  OR2X1 U9769 ( .A(n12685), .B(n10606), .Y(n13234) );
  NAND3X1 U9770 ( .A(n13225), .B(n11174), .C(n13234), .Y(n12686) );
  OAI21X1 U9771 ( .A(n12688), .B(n12687), .C(n12686), .Y(
        \lamb/scale_ls1/genblk1[1].mult/added[2] ) );
  AND2X1 U9772 ( .A(n13841), .B(\lamb/scale_ls1/genblk1[1].mult/added[2] ), 
        .Y(\lamb/scale_bs3/genblk1[1].mult/logA[2] ) );
  OAI21X1 U9773 ( .A(n10816), .B(n12690), .C(n10492), .Y(n12694) );
  NAND2X1 U9774 ( .A(n10816), .B(n12690), .Y(n12693) );
  AOI21X1 U9775 ( .A(n10817), .B(n12691), .C(n10549), .Y(n12692) );
  AOI21X1 U9776 ( .A(n12694), .B(n12693), .C(n12692), .Y(
        \lamb/scale_ts2/genblk1[2].mult/logA[2] ) );
  INVX1 U9777 ( .A(n13317), .Y(n13327) );
  AOI21X1 U9778 ( .A(n13225), .B(n12695), .C(n13327), .Y(n13246) );
  INVX1 U9779 ( .A(n13246), .Y(n13248) );
  AOI21X1 U9780 ( .A(n11227), .B(n13248), .C(n13857), .Y(n13132) );
  AOI22X1 U9781 ( .A(n13235), .B(n12696), .C(n13224), .D(n13324), .Y(n13243)
         );
  AOI22X1 U9782 ( .A(n12698), .B(n10828), .C(n13846), .D(n10591), .Y(n12708)
         );
  AOI21X1 U9783 ( .A(n13231), .B(n12699), .C(n13325), .Y(n13242) );
  OAI21X1 U9784 ( .A(n11169), .B(n13841), .C(n13848), .Y(n12705) );
  NAND2X1 U9785 ( .A(n12708), .B(n12705), .Y(n13129) );
  NAND2X1 U9786 ( .A(n13326), .B(n12700), .Y(n12703) );
  INVX1 U9787 ( .A(n12703), .Y(n13251) );
  OAI21X1 U9788 ( .A(n13841), .B(n13251), .C(n13855), .Y(n13131) );
  INVX1 U9789 ( .A(n13131), .Y(n13136) );
  INVX1 U9790 ( .A(n12705), .Y(n12706) );
  NAND2X1 U9791 ( .A(n13129), .B(n11015), .Y(n13128) );
  AOI22X1 U9792 ( .A(n13136), .B(n11015), .C(n13128), .D(n13131), .Y(n12702)
         );
  NAND2X1 U9793 ( .A(n10453), .B(n10579), .Y(n12704) );
  AOI22X1 U9794 ( .A(n13251), .B(n10827), .C(n10396), .D(n12704), .Y(
        \lamb/scale_ls2/genblk1[0].mult/logB[1] ) );
  NAND2X1 U9795 ( .A(n10594), .B(n12705), .Y(n12709) );
  OAI21X1 U9796 ( .A(n10824), .B(n12706), .C(n13131), .Y(n12707) );
  MUX2X1 U9797 ( .B(n10579), .A(n10828), .S(n10453), .Y(n12711) );
  AOI21X1 U9798 ( .A(n13251), .B(n10396), .C(n12711), .Y(
        \lamb/scale_ls2/genblk1[0].mult/logB[2] ) );
  AOI22X1 U9799 ( .A(n12715), .B(n12714), .C(n12954), .D(n12713), .Y(n12716)
         );
  OAI21X1 U9800 ( .A(n12717), .B(n11165), .C(n12716), .Y(n12718) );
  INVX1 U9801 ( .A(n12718), .Y(\forney/m0/logB [2]) );
  INVX1 U9802 ( .A(n13061), .Y(n13060) );
  INVX1 U9803 ( .A(n12719), .Y(n13052) );
  AOI21X1 U9804 ( .A(n13061), .B(n12720), .C(n13052), .Y(n12721) );
  MUX2X1 U9805 ( .B(n10651), .A(n13053), .S(n12721), .Y(n12722) );
  AOI21X1 U9806 ( .A(n13060), .B(n13064), .C(n12722), .Y(
        \lamb/scale_ds3/genblk1[3].mult/logA[2] ) );
  INVX1 U9807 ( .A(n13924), .Y(n12723) );
  NAND2X1 U9808 ( .A(n11119), .B(n10803), .Y(n13363) );
  NAND2X1 U9809 ( .A(n10600), .B(n13363), .Y(n13932) );
  AND2X1 U9810 ( .A(n12725), .B(n13932), .Y(n13364) );
  AOI21X1 U9811 ( .A(n11134), .B(n10803), .C(n13364), .Y(n12726) );
  INVX1 U9812 ( .A(n12726), .Y(\lamb/scale_ds1/genblk1[1].mult/logA[0] ) );
  INVX1 U9813 ( .A(\lamb/scale_ts1/genblk1[0].mult/added[1] ), .Y(n12745) );
  NAND2X1 U9814 ( .A(\lamb/scale_ts1/genblk1[0].mult/added[2] ), .B(n12745), 
        .Y(n12736) );
  INVX1 U9815 ( .A(n12736), .Y(n12732) );
  INVX1 U9816 ( .A(\add_x_145/n1 ), .Y(n12728) );
  INVX1 U9817 ( .A(\lamb/scale_ts1/genblk1[0].mult/added[3] ), .Y(n12735) );
  OR2X1 U9818 ( .A(\add_x_145/n1 ), .B(
        \lamb/scale_ts1/genblk1[0].mult/added[4] ), .Y(n12734) );
  NAND2X1 U9819 ( .A(\lamb/scale_ts1/genblk1[0].mult/added[4] ), .B(n12735), 
        .Y(n12727) );
  AOI22X1 U9820 ( .A(n12728), .B(n12735), .C(n12734), .D(n12727), .Y(n12754)
         );
  NAND2X1 U9821 ( .A(n12735), .B(n10513), .Y(n12730) );
  AND2X1 U9822 ( .A(\lamb/scale_ts1/genblk1[0].mult/added[3] ), .B(n12734), 
        .Y(n12741) );
  OAI21X1 U9823 ( .A(n12741), .B(\lamb/scale_ts1/genblk1[0].mult/added[2] ), 
        .C(\lamb/scale_ts1/genblk1[0].mult/added[1] ), .Y(n12729) );
  AOI21X1 U9824 ( .A(\lamb/scale_ts1/genblk1[0].mult/added[2] ), .B(n12730), 
        .C(n12729), .Y(n12731) );
  AOI21X1 U9825 ( .A(n12732), .B(n10784), .C(n12731), .Y(n12757) );
  NOR3X1 U9826 ( .A(\lamb/scale_ts1/genblk1[0].mult/added[3] ), .B(
        \add_x_145/n1 ), .C(\lamb/scale_ts1/genblk1[0].mult/added[4] ), .Y(
        n12742) );
  AOI21X1 U9827 ( .A(\lamb/scale_ts1/genblk1[0].mult/added[1] ), .B(n12742), 
        .C(n10784), .Y(n12733) );
  INVX1 U9828 ( .A(n12733), .Y(n12738) );
  NAND3X1 U9829 ( .A(\lamb/scale_ts1/genblk1[0].mult/added[3] ), .B(
        \add_x_145/n1 ), .C(\lamb/scale_ts1/genblk1[0].mult/added[4] ), .Y(
        n12739) );
  NAND3X1 U9830 ( .A(n12735), .B(n12734), .C(n10513), .Y(n12749) );
  AOI21X1 U9831 ( .A(n10751), .B(n12738), .C(n10912), .Y(n13210) );
  NAND2X1 U9832 ( .A(n12757), .B(n13210), .Y(n13209) );
  INVX1 U9833 ( .A(n13209), .Y(n13915) );
  INVX1 U9834 ( .A(n12742), .Y(n12744) );
  NAND3X1 U9835 ( .A(n12755), .B(n12744), .C(
        \lamb/scale_ts1/genblk1[0].mult/added[2] ), .Y(n12743) );
  OAI21X1 U9836 ( .A(\lamb/scale_ts1/genblk1[0].mult/added[2] ), .B(n10916), 
        .C(n12743), .Y(n12752) );
  OAI21X1 U9837 ( .A(n10751), .B(n10916), .C(n12744), .Y(n12748) );
  AOI21X1 U9838 ( .A(\lamb/scale_ts1/genblk1[0].mult/added[1] ), .B(n10784), 
        .C(n12748), .Y(n12747) );
  NAND2X1 U9839 ( .A(n12745), .B(n10916), .Y(n12746) );
  NAND2X1 U9840 ( .A(n13218), .B(n13917), .Y(n12759) );
  INVX1 U9841 ( .A(n12748), .Y(n12750) );
  AOI22X1 U9842 ( .A(\lamb/scale_ts1/genblk1[0].mult/added[1] ), .B(n12750), 
        .C(n10915), .D(n10751), .Y(n12751) );
  INVX1 U9843 ( .A(n13217), .Y(n13922) );
  OR2X1 U9844 ( .A(n10646), .B(n12759), .Y(n13219) );
  INVX1 U9845 ( .A(n13219), .Y(n12758) );
  AOI22X1 U9846 ( .A(\lamb/scale_ts1/genblk1[0].mult/added[1] ), .B(n10915), 
        .C(n12753), .D(n10784), .Y(n12756) );
  NAND3X1 U9847 ( .A(n12757), .B(n12756), .C(n12755), .Y(n13214) );
  INVX1 U9848 ( .A(n13214), .Y(n13914) );
  NOR2X1 U9849 ( .A(n11209), .B(n13914), .Y(n13216) );
  OAI21X1 U9850 ( .A(n13922), .B(n12758), .C(n13216), .Y(n13223) );
  OAI21X1 U9851 ( .A(n13915), .B(n12759), .C(n13223), .Y(
        \lamb/scale_ds2/genblk1[1].mult/logA[0] ) );
  AOI21X1 U9852 ( .A(n10528), .B(n13229), .C(n12760), .Y(n13228) );
  AOI21X1 U9853 ( .A(n13231), .B(n13314), .C(n13225), .Y(n12764) );
  MUX2X1 U9854 ( .B(n13229), .A(n13085), .S(n10749), .Y(n13241) );
  OAI21X1 U9855 ( .A(n13241), .B(n13083), .C(n10818), .Y(
        \lamb/scale_ls1/genblk1[1].mult/added[3] ) );
  INVX1 U9856 ( .A(\lamb/scale_ls1/genblk1[1].mult/added[3] ), .Y(n12763) );
  OAI21X1 U9857 ( .A(n11231), .B(n12763), .C(n13841), .Y(n13844) );
  NAND3X1 U9858 ( .A(\lamb/scale_ls2/genblk1[2].mult/added[1] ), .B(
        \lamb/scale_ls2/genblk1[2].mult/added[3] ), .C(
        \lamb/scale_ls2/genblk1[2].mult/added[2] ), .Y(n13107) );
  NOR2X1 U9859 ( .A(\lamb/scale_ls2/genblk1[2].mult/added[4] ), .B(
        \add_x_139/n1 ), .Y(n13108) );
  INVX1 U9860 ( .A(n13108), .Y(n12765) );
  NAND3X1 U9861 ( .A(n12765), .B(n11126), .C(n10673), .Y(n12766) );
  OAI21X1 U9862 ( .A(n11126), .B(n10673), .C(n12766), .Y(
        \lamb/scale_ls3/genblk1[2].mult/logA[3] ) );
  INVX1 U9863 ( .A(n12767), .Y(n13140) );
  AOI21X1 U9864 ( .A(n12768), .B(n11125), .C(n10820), .Y(n12769) );
  INVX1 U9865 ( .A(n12769), .Y(n12770) );
  NAND2X1 U9866 ( .A(n12858), .B(n11203), .Y(n12848) );
  NAND2X1 U9867 ( .A(n10699), .B(n10664), .Y(n13889) );
  INVX1 U9868 ( .A(n13889), .Y(n13897) );
  AOI21X1 U9869 ( .A(n11135), .B(n13897), .C(n10437), .Y(n13887) );
  AOI21X1 U9870 ( .A(n12771), .B(n10546), .C(n11210), .Y(n13905) );
  NOR2X1 U9871 ( .A(n13905), .B(n11172), .Y(n12774) );
  NAND2X1 U9872 ( .A(n12774), .B(n12772), .Y(n12773) );
  AOI21X1 U9873 ( .A(n10480), .B(n12773), .C(n10442), .Y(\forney/m0/logA [0])
         );
  OR2X1 U9874 ( .A(n12774), .B(n10582), .Y(n12776) );
  NAND2X1 U9875 ( .A(n10480), .B(\forney/m0/logA [3]), .Y(n12775) );
  OAI21X1 U9876 ( .A(n12776), .B(n11198), .C(n12775), .Y(\forney/m0/logA [2])
         );
  OR2X1 U9877 ( .A(\add_x_85/n1 ), .B(\forney/pe1/mult0/added [4]), .Y(n12892)
         );
  INVX1 U9878 ( .A(n12892), .Y(n12876) );
  INVX1 U9879 ( .A(\forney/pe1/mult0/added [3]), .Y(n12877) );
  INVX1 U9880 ( .A(\forney/pe1/mult0/added [1]), .Y(n12898) );
  NAND2X1 U9881 ( .A(n12881), .B(\forney/pe1/mult0/added [3]), .Y(n12777) );
  MUX2X1 U9882 ( .B(\forney/pe1/mult0/added [1]), .A(n12898), .S(n12777), .Y(
        n12778) );
  AOI22X1 U9883 ( .A(n12876), .B(n12877), .C(\forney/pe1/mult0/added [2]), .D(
        n12778), .Y(n12872) );
  NAND3X1 U9884 ( .A(n12779), .B(\forney/pe1/mult0/added [3]), .C(n12892), .Y(
        n12883) );
  NAND2X1 U9885 ( .A(n12876), .B(n12877), .Y(n12780) );
  NAND3X1 U9886 ( .A(\forney/pe1/mult0/added [2]), .B(n10435), .C(n12780), .Y(
        n12784) );
  AOI21X1 U9887 ( .A(n12881), .B(\forney/pe1/mult0/added [3]), .C(
        \forney/pe1/mult0/added [1]), .Y(n12782) );
  OAI21X1 U9888 ( .A(n12892), .B(n12877), .C(n11207), .Y(n12896) );
  INVX1 U9889 ( .A(n12896), .Y(n12781) );
  INVX1 U9890 ( .A(\forney/pe1/mult0/added [2]), .Y(n12893) );
  OAI21X1 U9891 ( .A(n12782), .B(n12781), .C(n12893), .Y(n12783) );
  NAND2X1 U9892 ( .A(n12784), .B(n12783), .Y(n12871) );
  INVX1 U9893 ( .A(n12871), .Y(n12785) );
  AOI21X1 U9894 ( .A(n11055), .B(\forney/pe1/mult0/added [1]), .C(n12785), .Y(
        n12843) );
  AND2X1 U9895 ( .A(n12892), .B(n12877), .Y(n12882) );
  NAND3X1 U9896 ( .A(n12882), .B(n12898), .C(n11207), .Y(n12890) );
  OR2X1 U9897 ( .A(n12804), .B(n13695), .Y(n12823) );
  AND2X1 U9898 ( .A(n13903), .B(n12823), .Y(n13901) );
  INVX1 U9899 ( .A(n13586), .Y(n12826) );
  NAND2X1 U9900 ( .A(n13891), .B(n13486), .Y(n12824) );
  NAND2X1 U9901 ( .A(n11210), .B(n12824), .Y(n13592) );
  INVX1 U9902 ( .A(n13592), .Y(n13694) );
  NAND2X1 U9903 ( .A(n10680), .B(n12809), .Y(n13692) );
  INVX1 U9904 ( .A(n13692), .Y(n12937) );
  AOI21X1 U9905 ( .A(n12858), .B(n10699), .C(n12937), .Y(n12788) );
  OAI21X1 U9906 ( .A(n12787), .B(n12788), .C(n12807), .Y(n12792) );
  INVX1 U9907 ( .A(n12824), .Y(n13908) );
  OAI21X1 U9908 ( .A(n13908), .B(n12790), .C(n12789), .Y(n12791) );
  AOI22X1 U9909 ( .A(n13694), .B(n12793), .C(n12792), .D(n12791), .Y(n12794)
         );
  AOI21X1 U9910 ( .A(n12826), .B(n12833), .C(n10910), .Y(n12798) );
  OR2X1 U9911 ( .A(n13488), .B(n12803), .Y(n13596) );
  OAI21X1 U9912 ( .A(n12795), .B(n13488), .C(n13596), .Y(n12796) );
  INVX1 U9913 ( .A(n12796), .Y(n12948) );
  AND2X1 U9914 ( .A(n10570), .B(n12948), .Y(n13697) );
  AOI22X1 U9915 ( .A(n13893), .B(n12798), .C(n13697), .D(n12797), .Y(n12802)
         );
  NAND2X1 U9916 ( .A(n10442), .B(n12799), .Y(n12801) );
  OAI21X1 U9917 ( .A(n10992), .B(n12802), .C(n12801), .Y(n12984) );
  INVX1 U9918 ( .A(n12984), .Y(n12989) );
  NAND2X1 U9919 ( .A(n13695), .B(n10477), .Y(n13579) );
  INVX1 U9920 ( .A(n13579), .Y(n12932) );
  NAND2X1 U9921 ( .A(n12804), .B(n12803), .Y(n12805) );
  HAX1 U9922 ( .A(n13488), .B(n12805), .YS(n12926) );
  AND2X1 U9923 ( .A(n12807), .B(n10546), .Y(n13589) );
  NOR2X1 U9924 ( .A(n13589), .B(n10680), .Y(n12808) );
  OAI21X1 U9925 ( .A(n11203), .B(n12809), .C(n12808), .Y(n12828) );
  NOR2X1 U9926 ( .A(n12829), .B(n12828), .Y(n12923) );
  NAND2X1 U9927 ( .A(n12826), .B(n12809), .Y(n12845) );
  AOI21X1 U9928 ( .A(n12845), .B(n12810), .C(n12858), .Y(n12811) );
  OR2X1 U9929 ( .A(n12923), .B(n12811), .Y(n12814) );
  INVX1 U9930 ( .A(n12812), .Y(n12813) );
  AOI22X1 U9931 ( .A(n13888), .B(n12814), .C(n13694), .D(n12813), .Y(n12817)
         );
  NAND3X1 U9932 ( .A(n13896), .B(n10798), .C(n10409), .Y(n12816) );
  NAND3X1 U9933 ( .A(n13582), .B(n12817), .C(n12816), .Y(n12818) );
  OAI21X1 U9934 ( .A(n12821), .B(n12926), .C(n12818), .Y(n12819) );
  OAI21X1 U9935 ( .A(n12821), .B(n10384), .C(n10873), .Y(n12992) );
  INVX1 U9936 ( .A(n12992), .Y(n12981) );
  OR2X1 U9937 ( .A(n12822), .B(n13903), .Y(n12930) );
  NOR2X1 U9938 ( .A(n13489), .B(n13888), .Y(n12825) );
  NOR2X1 U9939 ( .A(n11049), .B(n12825), .Y(n13601) );
  NAND3X1 U9940 ( .A(n12829), .B(n11129), .C(n12828), .Y(n12830) );
  NAND2X1 U9941 ( .A(n11161), .B(n12830), .Y(n12831) );
  OAI21X1 U9942 ( .A(n12832), .B(n11129), .C(n12831), .Y(n12835) );
  NOR3X1 U9943 ( .A(n12835), .B(n10833), .C(n10671), .Y(n12836) );
  AOI21X1 U9944 ( .A(n10833), .B(n12837), .C(n12836), .Y(n12838) );
  INVX1 U9945 ( .A(n12838), .Y(n12839) );
  AOI21X1 U9946 ( .A(n13601), .B(n12839), .C(n10564), .Y(n12840) );
  AOI21X1 U9947 ( .A(n10612), .B(n10698), .C(n12840), .Y(n12977) );
  AOI21X1 U9948 ( .A(n11084), .B(n10725), .C(n12842), .Y(n12903) );
  INVX1 U9949 ( .A(n10426), .Y(n12870) );
  AOI21X1 U9950 ( .A(n12843), .B(n12890), .C(n12870), .Y(n12869) );
  AOI22X1 U9951 ( .A(n10727), .B(n10564), .C(n11210), .D(n10798), .Y(n12866)
         );
  NAND2X1 U9952 ( .A(n12845), .B(n11195), .Y(n12846) );
  NOR3X1 U9953 ( .A(n11049), .B(n10753), .C(n12846), .Y(n12865) );
  INVX1 U9954 ( .A(n12848), .Y(n13591) );
  NAND2X1 U9955 ( .A(n10447), .B(n11161), .Y(n12851) );
  OAI21X1 U9956 ( .A(n12853), .B(n12852), .C(n12851), .Y(n12854) );
  AOI21X1 U9957 ( .A(n13591), .B(n12855), .C(n12854), .Y(n12942) );
  OAI21X1 U9958 ( .A(n11192), .B(n12857), .C(n12856), .Y(n12860) );
  NAND2X1 U9959 ( .A(n11192), .B(n12857), .Y(n12859) );
  NAND3X1 U9960 ( .A(n11025), .B(n12860), .C(n12859), .Y(n12861) );
  AOI21X1 U9961 ( .A(n12863), .B(n12862), .C(n12861), .Y(n12864) );
  HAX1 U9962 ( .A(n12869), .B(n10968), .YS(n13490) );
  INVX1 U9963 ( .A(n13490), .Y(n12912) );
  AOI21X1 U9964 ( .A(n11055), .B(n12871), .C(n12870), .Y(n12875) );
  NAND2X1 U9965 ( .A(n12873), .B(n12905), .Y(n12874) );
  HAX1 U9966 ( .A(n12875), .B(n12874), .YS(n13492) );
  AOI22X1 U9967 ( .A(n12912), .B(n13492), .C(n10854), .D(n13490), .Y(n12919)
         );
  AOI22X1 U9968 ( .A(\forney/pe1/mult0/added [3]), .B(n12876), .C(n12881), .D(
        n12877), .Y(n12891) );
  NAND3X1 U9969 ( .A(n12892), .B(n12893), .C(\forney/pe1/mult0/added [3]), .Y(
        n12897) );
  NAND3X1 U9970 ( .A(n11207), .B(n12877), .C(\forney/pe1/mult0/added [2]), .Y(
        n12878) );
  AOI21X1 U9971 ( .A(n10383), .B(n12878), .C(n12898), .Y(n12879) );
  INVX1 U9972 ( .A(n12879), .Y(n12901) );
  OAI21X1 U9973 ( .A(n12893), .B(n12891), .C(n12901), .Y(n12880) );
  INVX1 U9974 ( .A(n12880), .Y(n12885) );
  NAND3X1 U9975 ( .A(\forney/pe1/mult0/added [1]), .B(n12882), .C(n11207), .Y(
        n12884) );
  NAND3X1 U9976 ( .A(n12885), .B(n12884), .C(n10435), .Y(n12886) );
  NAND2X1 U9977 ( .A(n10426), .B(n12886), .Y(n12889) );
  NAND2X1 U9978 ( .A(n12887), .B(n12905), .Y(n12888) );
  HAX1 U9979 ( .A(n12889), .B(n12888), .YS(n12911) );
  INVX1 U9980 ( .A(n12911), .Y(n12917) );
  INVX1 U9981 ( .A(n12890), .Y(n12895) );
  OAI21X1 U9982 ( .A(n12898), .B(n12892), .C(n12891), .Y(n12894) );
  AOI22X1 U9983 ( .A(\forney/pe1/mult0/added [2]), .B(n12895), .C(n12894), .D(
        n12893), .Y(n12900) );
  NAND3X1 U9984 ( .A(n12898), .B(n10383), .C(n12896), .Y(n12899) );
  NAND2X1 U9985 ( .A(n10426), .B(n12902), .Y(n12907) );
  NAND2X1 U9986 ( .A(n12905), .B(n12904), .Y(n12906) );
  HAX1 U9987 ( .A(n12907), .B(n12906), .YS(n12916) );
  OAI21X1 U9988 ( .A(n10398), .B(n12917), .C(n11120), .Y(\forney/m1/logB [0])
         );
  NAND2X1 U9989 ( .A(n12912), .B(n11120), .Y(n12909) );
  OAI21X1 U9990 ( .A(n12917), .B(n13490), .C(n12916), .Y(n12908) );
  AOI22X1 U9991 ( .A(n12917), .B(n12909), .C(n13492), .D(n12908), .Y(
        \forney/m1/logB [1]) );
  AOI21X1 U9992 ( .A(n12912), .B(n12917), .C(n11120), .Y(n12915) );
  NAND2X1 U9993 ( .A(n12916), .B(n12911), .Y(n12920) );
  INVX1 U9994 ( .A(n12913), .Y(n12914) );
  NOR3X1 U9995 ( .A(n10439), .B(n12915), .C(n12914), .Y(\forney/m1/logB [2])
         );
  AND2X1 U9996 ( .A(n13490), .B(n10854), .Y(n12921) );
  OR2X1 U9997 ( .A(n12917), .B(n12916), .Y(n12918) );
  AOI22X1 U9998 ( .A(n12921), .B(n12920), .C(n10398), .D(n12918), .Y(
        \forney/m1/logB [3]) );
  AOI21X1 U9999 ( .A(n12922), .B(n10691), .C(n12923), .Y(n13575) );
  NOR2X1 U10000 ( .A(n11210), .B(n10671), .Y(n12924) );
  AOI22X1 U10001 ( .A(n13694), .B(n11060), .C(n13575), .D(n12924), .Y(n12928)
         );
  INVX1 U10002 ( .A(n12926), .Y(n13580) );
  AOI22X1 U10003 ( .A(n13582), .B(n12928), .C(n13580), .D(n10404), .Y(n12933)
         );
  AND2X1 U10004 ( .A(n12930), .B(n10582), .Y(n12931) );
  AOI22X1 U10005 ( .A(n12933), .B(n12932), .C(n12931), .D(n11198), .Y(
        \forney/m1/logA [1]) );
  NOR3X1 U10006 ( .A(n12937), .B(n12936), .C(n13750), .Y(n12939) );
  AOI22X1 U10007 ( .A(n13888), .B(n12939), .C(n12938), .D(n11210), .Y(n12940)
         );
  NAND3X1 U10008 ( .A(n11025), .B(n12941), .C(n12940), .Y(n12946) );
  INVX1 U10009 ( .A(n12943), .Y(n12945) );
  AOI22X1 U10010 ( .A(n13893), .B(n12946), .C(n12945), .D(n10570), .Y(n12947)
         );
  NAND3X1 U10011 ( .A(n12934), .B(n12948), .C(n12947), .Y(n12949) );
  OAI21X1 U10012 ( .A(n12950), .B(n13903), .C(n12949), .Y(n13912) );
  NOR2X1 U10013 ( .A(n10791), .B(n13912), .Y(\forney/m1/logA [3]) );
  OR2X1 U10014 ( .A(n12952), .B(n12951), .Y(n12957) );
  OAI21X1 U10015 ( .A(n12959), .B(n12955), .C(n12953), .Y(\forney/m0/logB [0])
         );
  INVX1 U10016 ( .A(n12954), .Y(n12960) );
  NAND2X1 U10017 ( .A(n11165), .B(n12955), .Y(n13480) );
  OAI21X1 U10018 ( .A(n12957), .B(n12960), .C(n13480), .Y(n12958) );
  AOI21X1 U10019 ( .A(n12960), .B(n12959), .C(n12958), .Y(\forney/m0/logB [3])
         );
  AOI21X1 U10020 ( .A(n12922), .B(n12963), .C(n10671), .Y(n12965) );
  AOI22X1 U10021 ( .A(n13486), .B(n12961), .C(n12965), .D(n12964), .Y(n12969)
         );
  OAI21X1 U10022 ( .A(n13896), .B(n12966), .C(n13488), .Y(n12967) );
  AOI22X1 U10023 ( .A(n11135), .B(n12969), .C(n12968), .D(n12967), .Y(n12972)
         );
  AOI22X1 U10024 ( .A(n13602), .B(n12972), .C(n10698), .D(n12971), .Y(n12973)
         );
  AOI21X1 U10025 ( .A(n13487), .B(n12974), .C(n12973), .Y(n12979) );
  INVX1 U10026 ( .A(n10725), .Y(n12983) );
  INVX1 U10027 ( .A(n10567), .Y(n12975) );
  NAND2X1 U10028 ( .A(n12981), .B(n12975), .Y(n12982) );
  OAI21X1 U10029 ( .A(n12976), .B(n12984), .C(n12982), .Y(
        \forney/pe1/mult0/logB [0]) );
  OAI21X1 U10030 ( .A(n10725), .B(n12984), .C(n12981), .Y(n12978) );
  AOI22X1 U10031 ( .A(n12981), .B(n12980), .C(n10567), .D(n12978), .Y(
        \forney/pe1/mult0/logB [1]) );
  AOI21X1 U10032 ( .A(n12989), .B(n12981), .C(n11176), .Y(n12986) );
  AOI21X1 U10033 ( .A(n12984), .B(n12983), .C(n12982), .Y(n12985) );
  NOR3X1 U10034 ( .A(n11084), .B(n12986), .C(n12985), .Y(
        \forney/pe1/mult0/logB [2]) );
  OAI21X1 U10035 ( .A(n12992), .B(n12988), .C(n12989), .Y(n12991) );
  AOI22X1 U10036 ( .A(n12988), .B(n12992), .C(n12991), .D(n11176), .Y(
        \forney/pe1/mult0/logB [3]) );
  OAI21X1 U10037 ( .A(n12799), .B(n11164), .C(n12993), .Y(n12995) );
  AOI21X1 U10038 ( .A(n11163), .B(n12995), .C(n12994), .Y(
        \forney/pe0/mult0/logB [1]) );
  NAND2X1 U10039 ( .A(n12799), .B(n13003), .Y(n12996) );
  MUX2X1 U10040 ( .B(n12997), .A(n11163), .S(n12996), .Y(n13000) );
  NAND3X1 U10041 ( .A(n12998), .B(n10659), .C(n13001), .Y(n12999) );
  OAI21X1 U10042 ( .A(n13001), .B(n13000), .C(n12999), .Y(
        \forney/pe0/mult0/logB [2]) );
  AOI21X1 U10043 ( .A(n13004), .B(n11164), .C(n13002), .Y(n13007) );
  OAI21X1 U10044 ( .A(n13007), .B(n10576), .C(n10659), .Y(
        \forney/pe0/mult0/logB [3]) );
  INVX1 U10045 ( .A(n13013), .Y(n13020) );
  AOI21X1 U10046 ( .A(n13008), .B(n13020), .C(n13015), .Y(n13010) );
  OAI21X1 U10047 ( .A(n13011), .B(n13010), .C(n13009), .Y(n13012) );
  INVX1 U10048 ( .A(n13012), .Y(\forney/pe0/mult0/logA [1]) );
  OAI21X1 U10049 ( .A(n13015), .B(n13014), .C(n13013), .Y(n13017) );
  NAND2X1 U10050 ( .A(n13015), .B(n13014), .Y(n13016) );
  NAND3X1 U10051 ( .A(n13018), .B(n13017), .C(n13016), .Y(n13019) );
  AOI21X1 U10052 ( .A(n10750), .B(n13020), .C(n13019), .Y(
        \forney/pe0/mult0/logA [2]) );
  OAI21X1 U10053 ( .A(n13023), .B(n10812), .C(n13022), .Y(
        \lamb/scale_ts3/genblk1[3].mult/logA[0] ) );
  NAND2X1 U10054 ( .A(n13027), .B(n10813), .Y(n13033) );
  OAI21X1 U10055 ( .A(n10813), .B(n10743), .C(n13024), .Y(n13026) );
  OAI21X1 U10056 ( .A(n10813), .B(n13027), .C(n13026), .Y(n13029) );
  INVX1 U10057 ( .A(n13031), .Y(n13032) );
  AOI21X1 U10058 ( .A(n13034), .B(n13033), .C(n13032), .Y(
        \lamb/scale_ts3/genblk1[3].mult/logA[3] ) );
  INVX1 U10059 ( .A(n10733), .Y(n13047) );
  AOI22X1 U10060 ( .A(n10830), .B(n13047), .C(n10733), .D(n10829), .Y(n13051)
         );
  INVX1 U10061 ( .A(n10690), .Y(n13043) );
  OAI21X1 U10062 ( .A(n13051), .B(n13043), .C(n10658), .Y(
        \lamb/scale_ts3/genblk1[2].mult/logA[0] ) );
  NOR3X1 U10063 ( .A(n10830), .B(n13043), .C(n13047), .Y(n13035) );
  NOR3X1 U10064 ( .A(n13037), .B(n10431), .C(n13035), .Y(
        \lamb/scale_ts3/genblk1[2].mult/logA[1] ) );
  NAND2X1 U10065 ( .A(n13038), .B(n10690), .Y(n13048) );
  NAND2X1 U10066 ( .A(n10733), .B(n13048), .Y(n13040) );
  MUX2X1 U10067 ( .B(n10830), .A(n10658), .S(n13040), .Y(n13042) );
  AOI21X1 U10068 ( .A(n13044), .B(n13043), .C(n13042), .Y(
        \lamb/scale_ts3/genblk1[2].mult/logA[2] ) );
  NAND2X1 U10069 ( .A(n10690), .B(n13044), .Y(n13050) );
  AND2X1 U10070 ( .A(n13047), .B(n10830), .Y(n13049) );
  AOI22X1 U10071 ( .A(n13051), .B(n13050), .C(n13049), .D(n13048), .Y(
        \lamb/scale_ts3/genblk1[2].mult/logA[3] ) );
  OR2X1 U10072 ( .A(n13052), .B(n13053), .Y(n13062) );
  OAI21X1 U10073 ( .A(n13064), .B(n13055), .C(n10651), .Y(
        \lamb/scale_ds3/genblk1[3].mult/logA[0] ) );
  NOR3X1 U10074 ( .A(n13058), .B(n13057), .C(n10966), .Y(
        \lamb/scale_ds3/genblk1[3].mult/logA[1] ) );
  MUX2X1 U10075 ( .B(n13061), .A(n13060), .S(n11095), .Y(n13063) );
  OAI21X1 U10076 ( .A(n13064), .B(n13063), .C(n13062), .Y(
        \lamb/scale_ds3/genblk1[3].mult/logA[3] ) );
  INVX1 U10077 ( .A(n13072), .Y(n13069) );
  OAI21X1 U10078 ( .A(n10822), .B(n13066), .C(n10650), .Y(
        \lamb/scale_ds3/genblk1[2].mult/logA[0] ) );
  OAI21X1 U10079 ( .A(n10724), .B(n10822), .C(n13077), .Y(n13068) );
  AOI21X1 U10080 ( .A(n13069), .B(n13068), .C(n13067), .Y(
        \lamb/scale_ds3/genblk1[2].mult/logA[1] ) );
  INVX1 U10081 ( .A(n13077), .Y(n13075) );
  AOI21X1 U10082 ( .A(n13077), .B(n13081), .C(n10724), .Y(n13071) );
  MUX2X1 U10083 ( .B(n10650), .A(n13072), .S(n13071), .Y(n13074) );
  AOI21X1 U10084 ( .A(n13075), .B(n10822), .C(n13074), .Y(
        \lamb/scale_ds3/genblk1[2].mult/logA[2] ) );
  AOI21X1 U10085 ( .A(n13078), .B(n13077), .C(n13076), .Y(n13080) );
  OAI21X1 U10086 ( .A(n10822), .B(n13080), .C(n10996), .Y(
        \lamb/scale_ds3/genblk1[2].mult/logA[3] ) );
  OAI21X1 U10087 ( .A(\lamb/scale_ls1/genblk1[1].mult/added[3] ), .B(
        \lamb/scale_ls1/genblk1[1].mult/added[2] ), .C(n10376), .Y(n13082) );
  INVX1 U10088 ( .A(n13082), .Y(n13842) );
  AOI21X1 U10089 ( .A(n13842), .B(n13085), .C(n13083), .Y(n13084) );
  OAI21X1 U10090 ( .A(n13842), .B(n13085), .C(n10874), .Y(n13087) );
  AOI21X1 U10091 ( .A(n10818), .B(n13087), .C(n11227), .Y(
        \lamb/scale_bs3/genblk1[1].mult/logA[3] ) );
  AOI22X1 U10092 ( .A(n13097), .B(n13098), .C(n13092), .D(n13091), .Y(n13103)
         );
  OAI21X1 U10093 ( .A(n10399), .B(n13101), .C(n10486), .Y(
        \lamb/scale_bs3/genblk1[0].mult/logB[0] ) );
  NAND2X1 U10094 ( .A(n13092), .B(n10486), .Y(n13089) );
  OAI21X1 U10095 ( .A(n13101), .B(n13098), .C(n13100), .Y(n13088) );
  AOI22X1 U10096 ( .A(n13101), .B(n13089), .C(n13091), .D(n13088), .Y(
        \lamb/scale_bs3/genblk1[0].mult/logB[1] ) );
  AOI21X1 U10097 ( .A(n13092), .B(n13101), .C(n10486), .Y(n13095) );
  NAND2X1 U10098 ( .A(n13092), .B(n13091), .Y(n13093) );
  AOI21X1 U10099 ( .A(n13099), .B(n13100), .C(n13093), .Y(n13094) );
  NOR3X1 U10100 ( .A(n11076), .B(n13095), .C(n13094), .Y(
        \lamb/scale_bs3/genblk1[0].mult/logB[2] ) );
  AND2X1 U10101 ( .A(n13098), .B(n13097), .Y(n13105) );
  NAND2X1 U10102 ( .A(n13099), .B(n13100), .Y(n13104) );
  OR2X1 U10103 ( .A(n13101), .B(n13100), .Y(n13102) );
  AOI22X1 U10104 ( .A(n13105), .B(n13104), .C(n10399), .D(n13102), .Y(
        \lamb/scale_bs3/genblk1[0].mult/logB[3] ) );
  INVX1 U10105 ( .A(\lamb/scale_ls2/genblk1[2].mult/added[1] ), .Y(n13109) );
  AND2X1 U10106 ( .A(\lamb/scale_ls2/genblk1[2].mult/added[3] ), .B(n13106), 
        .Y(n13114) );
  NAND2X1 U10107 ( .A(\lamb/scale_ls2/genblk1[2].mult/added[2] ), .B(n13114), 
        .Y(n13110) );
  AOI21X1 U10108 ( .A(n13109), .B(n13110), .C(n11136), .Y(
        \lamb/scale_ls3/genblk1[2].mult/logA[0] ) );
  OAI21X1 U10109 ( .A(\lamb/scale_ls2/genblk1[2].mult/added[2] ), .B(n13114), 
        .C(n13110), .Y(n13111) );
  NOR2X1 U10110 ( .A(\lamb/scale_ls2/genblk1[2].mult/added[3] ), .B(n13106), 
        .Y(n13112) );
  NOR3X1 U10111 ( .A(n13114), .B(n11136), .C(n13112), .Y(
        \lamb/scale_ls3/genblk1[2].mult/logA[2] ) );
  AOI21X1 U10112 ( .A(n13122), .B(n13121), .C(n11138), .Y(n13125) );
  OAI21X1 U10113 ( .A(n10402), .B(n13116), .C(n13115), .Y(
        \lamb/scale_ls3/genblk1[1].mult/logA[0] ) );
  INVX1 U10114 ( .A(n13116), .Y(n13867) );
  NAND2X1 U10115 ( .A(n13119), .B(n13867), .Y(n13126) );
  OAI21X1 U10116 ( .A(n13867), .B(n13121), .C(n13117), .Y(n13118) );
  OAI21X1 U10117 ( .A(n13867), .B(n13119), .C(n13118), .Y(n13120) );
  AOI21X1 U10118 ( .A(n11138), .B(n13126), .C(n13120), .Y(
        \lamb/scale_ls3/genblk1[1].mult/logA[2] ) );
  AND2X1 U10119 ( .A(n13122), .B(n13121), .Y(n13127) );
  AOI22X1 U10120 ( .A(n13127), .B(n13126), .C(n10402), .D(n10943), .Y(
        \lamb/scale_ls3/genblk1[1].mult/logA[3] ) );
  INVX1 U10121 ( .A(n13128), .Y(n13130) );
  OAI21X1 U10122 ( .A(n10824), .B(n13130), .C(n10594), .Y(
        \lamb/scale_ls3/genblk1[0].mult/logB[0] ) );
  AND2X1 U10123 ( .A(n13131), .B(n13130), .Y(n13133) );
  MUX2X1 U10124 ( .B(n10594), .A(n13133), .S(n10824), .Y(n13135) );
  AOI21X1 U10125 ( .A(n13136), .B(n10838), .C(n13135), .Y(
        \lamb/scale_ls3/genblk1[0].mult/logB[2] ) );
  OAI21X1 U10126 ( .A(n10483), .B(n10820), .C(n13143), .Y(n13139) );
  AOI21X1 U10127 ( .A(n13140), .B(n13139), .C(n13138), .Y(
        \lamb/scale_ls3/genblk1[0].mult/logA[1] ) );
  NOR2X1 U10128 ( .A(n13141), .B(n11177), .Y(n13146) );
  AOI21X1 U10129 ( .A(n13143), .B(n10819), .C(n11125), .Y(n13145) );
  AOI22X1 U10130 ( .A(n10820), .B(n13143), .C(n11177), .D(n10819), .Y(n13144)
         );
  NOR3X1 U10131 ( .A(n13146), .B(n13145), .C(n13144), .Y(
        \lamb/scale_ls3/genblk1[0].mult/logA[2] ) );
  NOR2X1 U10132 ( .A(n13147), .B(n13146), .Y(n13149) );
  OAI21X1 U10133 ( .A(n10820), .B(n13149), .C(n11125), .Y(
        \lamb/scale_ls3/genblk1[0].mult/logA[3] ) );
  NAND2X1 U10134 ( .A(n13161), .B(n13158), .Y(n13153) );
  OAI21X1 U10135 ( .A(n13152), .B(n13151), .C(n13153), .Y(
        \lamb/scale_ts2/genblk1[3].mult/logA[0] ) );
  AOI21X1 U10136 ( .A(n13154), .B(n13153), .C(n13157), .Y(n13156) );
  INVX1 U10137 ( .A(n13156), .Y(n13166) );
  NAND2X1 U10138 ( .A(n13158), .B(n13157), .Y(n13170) );
  INVX1 U10139 ( .A(n13170), .Y(n13164) );
  OAI21X1 U10140 ( .A(n13161), .B(n13160), .C(n10995), .Y(n13162) );
  OAI21X1 U10141 ( .A(n13164), .B(n11031), .C(n13162), .Y(n13165) );
  OAI21X1 U10142 ( .A(n13167), .B(n13166), .C(n13165), .Y(
        \lamb/scale_ts2/genblk1[3].mult/logA[2] ) );
  INVX1 U10143 ( .A(n13168), .Y(n13171) );
  AOI21X1 U10144 ( .A(n13171), .B(n13170), .C(n13169), .Y(
        \lamb/scale_ts2/genblk1[3].mult/logA[3] ) );
  NOR3X1 U10145 ( .A(n10425), .B(n10432), .C(n11042), .Y(
        \lamb/scale_ts2/genblk1[2].mult/logA[1] ) );
  NAND2X1 U10146 ( .A(n10732), .B(n13868), .Y(n13174) );
  HAX1 U10147 ( .A(n10726), .B(n13174), .YS(n13177) );
  OAI21X1 U10148 ( .A(n10817), .B(n13177), .C(n10492), .Y(
        \lamb/scale_ts2/genblk1[2].mult/logA[3] ) );
  INVX1 U10149 ( .A(n10703), .Y(n13180) );
  NAND2X1 U10150 ( .A(n10800), .B(n10805), .Y(n13944) );
  NAND3X1 U10151 ( .A(n13180), .B(n10832), .C(n13944), .Y(n13182) );
  AOI21X1 U10152 ( .A(n11056), .B(n13182), .C(n13179), .Y(
        \lamb/scale_ts2/genblk1[1].mult/logA[1] ) );
  NAND2X1 U10153 ( .A(n13180), .B(n10832), .Y(n13181) );
  OAI21X1 U10154 ( .A(n10800), .B(n10804), .C(n13181), .Y(n13183) );
  NAND2X1 U10155 ( .A(n13183), .B(n13182), .Y(n13184) );
  OAI21X1 U10156 ( .A(n11056), .B(n10805), .C(n13184), .Y(
        \lamb/scale_ts2/genblk1[1].mult/logA[2] ) );
  MUX2X1 U10157 ( .B(n10805), .A(n10804), .S(n10495), .Y(n13189) );
  OAI21X1 U10158 ( .A(n10832), .B(n13189), .C(n13943), .Y(
        \lamb/scale_ts2/genblk1[1].mult/logA[3] ) );
  AOI22X1 U10159 ( .A(n13880), .B(n13191), .C(n13876), .D(n13877), .Y(n13197)
         );
  OAI21X1 U10160 ( .A(n10400), .B(n13879), .C(n11121), .Y(
        \lamb/scale_ds2/genblk1[3].mult/logA[0] ) );
  NAND2X1 U10161 ( .A(n13880), .B(n11121), .Y(n13192) );
  OAI21X1 U10162 ( .A(n13879), .B(n13877), .C(n13193), .Y(n13190) );
  AOI22X1 U10163 ( .A(n13879), .B(n13192), .C(n13191), .D(n13190), .Y(
        \lamb/scale_ds2/genblk1[3].mult/logA[1] ) );
  AND2X1 U10164 ( .A(n13877), .B(n13876), .Y(n13198) );
  NAND2X1 U10165 ( .A(n13193), .B(n13195), .Y(n13885) );
  NAND2X1 U10166 ( .A(n13195), .B(n13194), .Y(n13196) );
  AOI22X1 U10167 ( .A(n13198), .B(n13885), .C(n10400), .D(n13196), .Y(
        \lamb/scale_ds2/genblk1[3].mult/logA[3] ) );
  AOI21X1 U10168 ( .A(n13933), .B(n13935), .C(n11139), .Y(n13208) );
  OAI21X1 U10169 ( .A(n10381), .B(n13200), .C(n13199), .Y(
        \lamb/scale_ds2/genblk1[2].mult/logA[0] ) );
  OR2X1 U10170 ( .A(n13202), .B(n13201), .Y(n13203) );
  AOI21X1 U10171 ( .A(n11139), .B(n13934), .C(n13203), .Y(
        \lamb/scale_ds2/genblk1[2].mult/logA[1] ) );
  AOI22X1 U10172 ( .A(n10381), .B(n10403), .C(n10941), .D(n10407), .Y(
        \lamb/scale_ds2/genblk1[2].mult/logA[3] ) );
  NAND2X1 U10173 ( .A(n13917), .B(n13209), .Y(n13222) );
  INVX1 U10174 ( .A(n13917), .Y(n13212) );
  NAND2X1 U10175 ( .A(n13212), .B(n13210), .Y(n13211) );
  NAND2X1 U10176 ( .A(n13212), .B(n13915), .Y(n13213) );
  NAND3X1 U10177 ( .A(n13214), .B(n13217), .C(n13213), .Y(n13215) );
  AOI21X1 U10178 ( .A(n13918), .B(n13215), .C(n11209), .Y(
        \lamb/scale_ds2/genblk1[1].mult/logA[1] ) );
  NAND2X1 U10179 ( .A(n13915), .B(n13216), .Y(n13921) );
  OAI21X1 U10180 ( .A(n11209), .B(n13217), .C(n13921), .Y(n13220) );
  NAND2X1 U10181 ( .A(n13220), .B(n13219), .Y(n13221) );
  OAI21X1 U10182 ( .A(n13223), .B(n13222), .C(n13221), .Y(
        \lamb/scale_ds2/genblk1[1].mult/logA[3] ) );
  AND2X1 U10183 ( .A(n13231), .B(n13314), .Y(n13226) );
  NAND3X1 U10184 ( .A(n13226), .B(n10809), .C(n10826), .Y(n13227) );
  OAI21X1 U10185 ( .A(n10826), .B(n13228), .C(n13227), .Y(
        \lamb/scale_bs2/genblk1[0].mult/logA[1] ) );
  NAND2X1 U10186 ( .A(n13229), .B(n10818), .Y(n13237) );
  AOI21X1 U10187 ( .A(n10826), .B(n13231), .C(n11174), .Y(n13232) );
  INVX1 U10188 ( .A(n13232), .Y(n13233) );
  NAND3X1 U10189 ( .A(n10809), .B(n13234), .C(n13233), .Y(n13236) );
  AOI21X1 U10190 ( .A(n13237), .B(n10826), .C(n13236), .Y(
        \lamb/scale_bs2/genblk1[0].mult/logA[2] ) );
  OR2X1 U10191 ( .A(n10818), .B(n13235), .Y(n13239) );
  OAI21X1 U10192 ( .A(n13241), .B(n10826), .C(n13239), .Y(
        \lamb/scale_bs2/genblk1[0].mult/logA[3] ) );
  NAND2X1 U10193 ( .A(n10828), .B(n11169), .Y(n13247) );
  AND2X1 U10194 ( .A(n13249), .B(n13247), .Y(n13245) );
  OAI21X1 U10195 ( .A(n13246), .B(n13245), .C(n10579), .Y(
        \lamb/scale_ls2/genblk1[0].mult/logB[0] ) );
  INVX1 U10196 ( .A(n13247), .Y(n13252) );
  OAI21X1 U10197 ( .A(n13251), .B(n13252), .C(n13248), .Y(n13250) );
  AOI22X1 U10198 ( .A(n13252), .B(n13251), .C(n13250), .D(n13249), .Y(
        \lamb/scale_ls2/genblk1[0].mult/logB[3] ) );
  NAND2X1 U10199 ( .A(n13325), .B(n13317), .Y(n13322) );
  NAND2X1 U10200 ( .A(n13253), .B(n13322), .Y(n13254) );
  NAND3X1 U10201 ( .A(n13256), .B(n11124), .C(n13254), .Y(n13257) );
  OAI21X1 U10202 ( .A(n13259), .B(n10627), .C(n13257), .Y(
        \lamb/scale_ls2/genblk1[0].mult/logA[2] ) );
  AOI22X1 U10203 ( .A(n13273), .B(n13272), .C(n13267), .D(n13262), .Y(n13277)
         );
  OAI21X1 U10204 ( .A(n10401), .B(n10471), .C(n13260), .Y(
        \lamb/scale_ts1/genblk1[2].mult/logA[0] ) );
  NOR2X1 U10205 ( .A(n13262), .B(n13267), .Y(n13271) );
  NAND2X1 U10206 ( .A(n11020), .B(n13263), .Y(n13265) );
  AOI21X1 U10207 ( .A(n13274), .B(n13271), .C(n13265), .Y(
        \lamb/scale_ts1/genblk1[2].mult/logA[1] ) );
  OAI21X1 U10208 ( .A(n13267), .B(n13274), .C(n13266), .Y(n13268) );
  OAI21X1 U10209 ( .A(n13274), .B(n13269), .C(n13268), .Y(n13270) );
  AOI21X1 U10210 ( .A(n13271), .B(n11058), .C(n13270), .Y(
        \lamb/scale_ts1/genblk1[2].mult/logA[2] ) );
  NOR2X1 U10211 ( .A(n13273), .B(n13272), .Y(n13279) );
  NAND2X1 U10212 ( .A(n13275), .B(n13274), .Y(n13276) );
  AOI22X1 U10213 ( .A(n13279), .B(n11058), .C(n10401), .D(n13276), .Y(
        \lamb/scale_ts1/genblk1[2].mult/logA[3] ) );
  OAI21X1 U10214 ( .A(n11071), .B(n10796), .C(n10657), .Y(
        \lamb/scale_ts1/genblk1[1].mult/logA[0] ) );
  NOR3X1 U10215 ( .A(n11075), .B(n10796), .C(n10794), .Y(n13281) );
  NOR3X1 U10216 ( .A(n10424), .B(n10430), .C(n13281), .Y(
        \lamb/scale_ts1/genblk1[1].mult/logA[1] ) );
  NAND2X1 U10217 ( .A(n10808), .B(n10797), .Y(n13290) );
  NAND2X1 U10218 ( .A(n10795), .B(n13290), .Y(n13285) );
  MUX2X1 U10219 ( .B(n11075), .A(n10657), .S(n13285), .Y(n13287) );
  AOI21X1 U10220 ( .A(n10681), .B(n10796), .C(n13287), .Y(
        \lamb/scale_ts1/genblk1[1].mult/logA[2] ) );
  NAND2X1 U10221 ( .A(n10797), .B(n10681), .Y(n13292) );
  AND2X1 U10222 ( .A(n10794), .B(n11075), .Y(n13291) );
  AOI22X1 U10223 ( .A(n11071), .B(n13292), .C(n13291), .D(n13290), .Y(
        \lamb/scale_ts1/genblk1[1].mult/logA[3] ) );
  INVX1 U10224 ( .A(n13296), .Y(n13295) );
  AOI22X1 U10225 ( .A(msg[2]), .B(msg[25]), .C(n13723), .D(n13811), .Y(n13294)
         );
  MUX2X1 U10226 ( .B(n13296), .A(n13295), .S(n13294), .Y(n13297) );
  MUX2X1 U10227 ( .B(n13299), .A(n13298), .S(n13297), .Y(n13309) );
  MUX2X1 U10228 ( .B(n13300), .A(msg[59]), .S(msg[49]), .Y(n13301) );
  FAX1 U10229 ( .A(n13303), .B(n13302), .C(n13301), .YS(n13304) );
  MUX2X1 U10230 ( .B(n13306), .A(n13305), .S(n13304), .Y(n13307) );
  FAX1 U10231 ( .A(n13309), .B(n11150), .C(n13307), .YS(n13310) );
  FAX1 U10232 ( .A(n13312), .B(n13311), .C(n13310), .YS(n13313) );
  MUX2X1 U10233 ( .B(n13314), .A(n10674), .S(n13313), .Y(n13329) );
  NOR2X1 U10234 ( .A(n13326), .B(n13324), .Y(n13323) );
  OAI21X1 U10235 ( .A(n13317), .B(n13329), .C(n11219), .Y(
        \lamb/scale_ts1/genblk1[0].mult/logB[0] ) );
  NAND2X1 U10236 ( .A(n13325), .B(n11219), .Y(n13316) );
  INVX1 U10237 ( .A(n13326), .Y(n13318) );
  OAI21X1 U10238 ( .A(n13316), .B(n13317), .C(n13318), .Y(n13315) );
  AOI22X1 U10239 ( .A(n13317), .B(n13316), .C(n13315), .D(n13324), .Y(
        \lamb/scale_ts1/genblk1[0].mult/logB[1] ) );
  NAND3X1 U10240 ( .A(n13324), .B(n13325), .C(n10420), .Y(n13320) );
  NAND2X1 U10241 ( .A(n13320), .B(n10440), .Y(n13321) );
  NOR2X1 U10242 ( .A(n13325), .B(n13324), .Y(n13331) );
  NAND2X1 U10243 ( .A(n13327), .B(n13326), .Y(n13328) );
  AOI22X1 U10244 ( .A(n13331), .B(n10420), .C(n13329), .D(n13328), .Y(
        \lamb/scale_ts1/genblk1[0].mult/logB[3] ) );
  INVX1 U10245 ( .A(n13336), .Y(n13831) );
  NAND2X1 U10246 ( .A(n13333), .B(n11117), .Y(n13836) );
  NAND3X1 U10247 ( .A(n13831), .B(n13830), .C(n11137), .Y(n13335) );
  AOI21X1 U10248 ( .A(n13836), .B(n13335), .C(n13334), .Y(
        \lamb/scale_ds1/genblk1[3].mult/logA[1] ) );
  MUX2X1 U10249 ( .B(n13337), .A(n13837), .S(n10498), .Y(n13338) );
  OAI21X1 U10250 ( .A(n13830), .B(n13338), .C(n11117), .Y(
        \lamb/scale_ds1/genblk1[3].mult/logA[3] ) );
  INVX1 U10251 ( .A(n13348), .Y(n13874) );
  NOR2X1 U10252 ( .A(n13874), .B(n11118), .Y(n13339) );
  NOR3X1 U10253 ( .A(n13341), .B(n13340), .C(n13339), .Y(
        \lamb/scale_ds1/genblk1[2].mult/logA[1] ) );
  OAI21X1 U10254 ( .A(n13342), .B(n13348), .C(n11118), .Y(n13344) );
  AOI21X1 U10255 ( .A(n13350), .B(n13874), .C(n10626), .Y(n13343) );
  AOI21X1 U10256 ( .A(n11078), .B(n13344), .C(n13343), .Y(
        \lamb/scale_ds1/genblk1[2].mult/logA[2] ) );
  OAI21X1 U10257 ( .A(n13349), .B(n13350), .C(n11118), .Y(n13346) );
  INVX1 U10258 ( .A(n13346), .Y(n13875) );
  NAND2X1 U10259 ( .A(n13348), .B(n13347), .Y(n13353) );
  NOR2X1 U10260 ( .A(n13350), .B(n13349), .Y(n13352) );
  AOI22X1 U10261 ( .A(n13875), .B(n13353), .C(n13352), .D(n11078), .Y(
        \lamb/scale_ds1/genblk1[2].mult/logA[3] ) );
  AOI21X1 U10262 ( .A(n13354), .B(n13355), .C(n13925), .Y(n13360) );
  AOI21X1 U10263 ( .A(n13355), .B(n13925), .C(n10468), .Y(n13365) );
  OAI21X1 U10264 ( .A(n11119), .B(n10803), .C(n10474), .Y(n13357) );
  NAND2X1 U10265 ( .A(n13365), .B(n13357), .Y(n13358) );
  OAI21X1 U10266 ( .A(n13360), .B(n13359), .C(n13358), .Y(
        \lamb/scale_ds1/genblk1[1].mult/logA[1] ) );
  OAI21X1 U10267 ( .A(n11134), .B(n10474), .C(n10600), .Y(n13928) );
  AOI22X1 U10268 ( .A(n13365), .B(n13364), .C(n13363), .D(n13928), .Y(n13366)
         );
  INVX1 U10269 ( .A(n13366), .Y(\lamb/scale_ds1/genblk1[1].mult/logA[3] ) );
  OAI21X1 U10270 ( .A(n13826), .B(n13367), .C(n13370), .Y(n13369) );
  AOI21X1 U10271 ( .A(n13372), .B(n13369), .C(n13368), .Y(
        \lamb/scale_ts0/genblk1[1].mult/logA[1] ) );
  OAI21X1 U10272 ( .A(n13370), .B(n13377), .C(n10501), .Y(n13375) );
  NAND2X1 U10273 ( .A(n13370), .B(n13377), .Y(n13374) );
  OAI21X1 U10274 ( .A(n13372), .B(n13374), .C(n13376), .Y(n13373) );
  AOI21X1 U10275 ( .A(n13375), .B(n13374), .C(n13373), .Y(
        \lamb/scale_ts0/genblk1[1].mult/logA[2] ) );
  INVX1 U10276 ( .A(n13376), .Y(n13379) );
  OAI21X1 U10277 ( .A(n13379), .B(n13378), .C(n13377), .Y(n13380) );
  NAND2X1 U10278 ( .A(n10501), .B(n13380), .Y(
        \lamb/scale_ts0/genblk1[1].mult/logA[3] ) );
  NOR3X1 U10279 ( .A(n12682), .B(n11024), .C(n10630), .Y(n13383) );
  INVX1 U10280 ( .A(n13383), .Y(n13384) );
  OAI21X1 U10281 ( .A(n13385), .B(n13384), .C(n13602), .Y(n13751) );
  NOR2X1 U10282 ( .A(n10833), .B(n13751), .Y(n13386) );
  NAND2X1 U10283 ( .A(n13387), .B(n13386), .Y(valid) );
  AND2X1 U10284 ( .A(\forney/m0/added [4]), .B(\add_x_14/n1 ), .Y(n13392) );
  NOR2X1 U10285 ( .A(\forney/m0/added [3]), .B(n13392), .Y(n13390) );
  INVX1 U10286 ( .A(n13390), .Y(n13408) );
  OR2X1 U10287 ( .A(\forney/m0/added [4]), .B(\add_x_14/n1 ), .Y(n13389) );
  INVX1 U10288 ( .A(\forney/m0/added [2]), .Y(n13417) );
  MUX2X1 U10289 ( .B(n13408), .A(n11141), .S(n13417), .Y(n13388) );
  NAND2X1 U10290 ( .A(\forney/m0/added [1]), .B(n13388), .Y(n13421) );
  NAND2X1 U10291 ( .A(n13390), .B(n13389), .Y(n13396) );
  INVX1 U10292 ( .A(n13396), .Y(n13401) );
  INVX1 U10293 ( .A(n10382), .Y(n13397) );
  AOI22X1 U10294 ( .A(\forney/m0/added [1]), .B(n13401), .C(
        \forney/m0/added [2]), .D(n13397), .Y(n13394) );
  NOR3X1 U10295 ( .A(\forney/m0/added [1]), .B(n13392), .C(n11141), .Y(n13393)
         );
  INVX1 U10296 ( .A(n13393), .Y(n13395) );
  NOR3X1 U10297 ( .A(\forney/m0/added [3]), .B(\forney/m0/added [4]), .C(
        \add_x_14/n1 ), .Y(n13399) );
  INVX1 U10298 ( .A(n13399), .Y(n13415) );
  AOI21X1 U10299 ( .A(n13415), .B(n13395), .C(n13417), .Y(n13410) );
  NAND3X1 U10300 ( .A(\forney/m0/added [3]), .B(\forney/m0/added [4]), .C(
        \add_x_14/n1 ), .Y(n13405) );
  NAND2X1 U10301 ( .A(n13397), .B(\forney/m0/added [1]), .Y(n13398) );
  AOI21X1 U10302 ( .A(n13413), .B(n13398), .C(\forney/m0/added [2]), .Y(n13407) );
  INVX1 U10303 ( .A(n10991), .Y(n13403) );
  INVX1 U10304 ( .A(\forney/m0/added [1]), .Y(n13419) );
  NOR2X1 U10305 ( .A(n13419), .B(n13417), .Y(n13400) );
  AOI21X1 U10306 ( .A(n13400), .B(n10644), .C(n13399), .Y(n13404) );
  AOI22X1 U10307 ( .A(\forney/m0/added [1]), .B(n11014), .C(n13401), .D(n13419), .Y(n13402) );
  NAND2X1 U10308 ( .A(n13403), .B(n13402), .Y(n13412) );
  NOR2X1 U10309 ( .A(n13410), .B(n13412), .Y(n13424) );
  OAI21X1 U10310 ( .A(\forney/m0/added [1]), .B(n10644), .C(n11014), .Y(n13406) );
  AOI21X1 U10311 ( .A(n13408), .B(n10991), .C(n13406), .Y(n13409) );
  INVX1 U10312 ( .A(n13409), .Y(n13411) );
  NAND2X1 U10313 ( .A(n10534), .B(n10445), .Y(n13422) );
  OAI21X1 U10314 ( .A(n13413), .B(n13417), .C(n10382), .Y(n13418) );
  OAI21X1 U10315 ( .A(n13419), .B(n13415), .C(n10382), .Y(n13416) );
  AOI22X1 U10316 ( .A(n13419), .B(n13418), .C(n13417), .D(n13416), .Y(n13420)
         );
  NOR2X1 U10317 ( .A(n11202), .B(n13450), .Y(n13448) );
  AOI21X1 U10318 ( .A(n13443), .B(n13422), .C(n13448), .Y(n13469) );
  NOR2X1 U10319 ( .A(n13437), .B(n13478), .Y(n13435) );
  AOI21X1 U10320 ( .A(n13436), .B(n11196), .C(n13435), .Y(n13423) );
  INVX1 U10321 ( .A(n13423), .Y(n13549) );
  OAI21X1 U10322 ( .A(n11202), .B(n13450), .C(n10662), .Y(n13425) );
  AOI22X1 U10323 ( .A(n13450), .B(n11202), .C(n13425), .D(n10438), .Y(n13472)
         );
  AND2X1 U10324 ( .A(n13427), .B(n13426), .Y(n13428) );
  AOI21X1 U10325 ( .A(n13429), .B(n13436), .C(n13428), .Y(n13530) );
  NAND2X1 U10326 ( .A(n13458), .B(n13439), .Y(n13434) );
  INVX1 U10327 ( .A(n13430), .Y(n13432) );
  OAI21X1 U10328 ( .A(n13432), .B(n13431), .C(n10585), .Y(n13433) );
  AOI21X1 U10329 ( .A(n13435), .B(n13434), .C(n13433), .Y(n13538) );
  AND2X1 U10330 ( .A(n13437), .B(n13436), .Y(n13441) );
  OAI21X1 U10331 ( .A(n13439), .B(n13441), .C(n13438), .Y(n13440) );
  OAI21X1 U10332 ( .A(n11196), .B(n13441), .C(n13440), .Y(n13535) );
  INVX1 U10333 ( .A(n13443), .Y(n13447) );
  HAX1 U10334 ( .A(n10534), .B(n13450), .YS(n13446) );
  OAI21X1 U10335 ( .A(n13447), .B(n13446), .C(n10445), .Y(n13476) );
  NAND2X1 U10336 ( .A(n13535), .B(n13476), .Y(n13455) );
  NAND2X1 U10337 ( .A(n11162), .B(n13455), .Y(n13462) );
  INVX1 U10338 ( .A(n13462), .Y(n13456) );
  INVX1 U10339 ( .A(n13448), .Y(n13453) );
  AOI22X1 U10340 ( .A(n10662), .B(n11202), .C(n13450), .D(n10438), .Y(n13452)
         );
  OAI21X1 U10341 ( .A(n10662), .B(n13453), .C(n13452), .Y(n13465) );
  OAI21X1 U10342 ( .A(n13456), .B(n13465), .C(n13463), .Y(n13457) );
  OR2X1 U10343 ( .A(n13457), .B(n10456), .Y(n13470) );
  OAI21X1 U10344 ( .A(n10697), .B(n13471), .C(n13470), .Y(n13460) );
  OR2X1 U10345 ( .A(n13549), .B(n13460), .Y(n13468) );
  AOI21X1 U10346 ( .A(n13549), .B(n13460), .C(n11158), .Y(n13466) );
  NAND2X1 U10347 ( .A(n13468), .B(n13466), .Y(n13461) );
  HAX1 U10348 ( .A(n10640), .B(n13461), .YS(n13626) );
  INVX1 U10349 ( .A(n13626), .Y(n13605) );
  NAND3X1 U10350 ( .A(n13547), .B(n13463), .C(n13462), .Y(n13464) );
  HAX1 U10351 ( .A(n13465), .B(n13464), .YS(n13628) );
  INVX1 U10352 ( .A(n13628), .Y(n13609) );
  AND2X1 U10353 ( .A(n13605), .B(n10811), .Y(n13475) );
  INVX1 U10354 ( .A(n13466), .Y(n13467) );
  AOI21X1 U10355 ( .A(n10640), .B(n13468), .C(n13467), .Y(n13634) );
  NAND3X1 U10356 ( .A(n13547), .B(n10998), .C(n13470), .Y(n13473) );
  XNOR2X1 U10357 ( .A(n13473), .B(n10697), .Y(n13627) );
  NAND3X1 U10358 ( .A(n11208), .B(n13627), .C(n10811), .Y(n13474) );
  OAI21X1 U10359 ( .A(n13475), .B(n11208), .C(n13474), .Y(n13482) );
  INVX1 U10360 ( .A(n13476), .Y(n13477) );
  HAX1 U10361 ( .A(n13477), .B(n10655), .YS(n13631) );
  OAI21X1 U10362 ( .A(n11208), .B(n13627), .C(n10811), .Y(n13651) );
  NAND2X1 U10363 ( .A(n11158), .B(n13478), .Y(n13494) );
  OAI21X1 U10364 ( .A(n13480), .B(n13479), .C(n13494), .Y(n13650) );
  AOI21X1 U10365 ( .A(n13651), .B(n13631), .C(n13650), .Y(n13481) );
  OAI21X1 U10366 ( .A(n13482), .B(n13631), .C(n13481), .Y(n13702) );
  OAI21X1 U10367 ( .A(n10691), .B(n10573), .C(n10699), .Y(n13576) );
  OAI21X1 U10368 ( .A(n13486), .B(n13576), .C(n13896), .Y(n13684) );
  AOI21X1 U10369 ( .A(n13488), .B(n13684), .C(n13487), .Y(n13574) );
  AOI21X1 U10370 ( .A(n10664), .B(n13888), .C(n10727), .Y(n13667) );
  INVX1 U10371 ( .A(n13667), .Y(n13753) );
  NAND3X1 U10372 ( .A(n13492), .B(n10439), .C(n13490), .Y(n13493) );
  INVX1 U10373 ( .A(\forney/m1/added [3]), .Y(n13504) );
  AOI22X1 U10374 ( .A(\forney/m1/added [3]), .B(n11197), .C(n13496), .D(n13504), .Y(n13516) );
  INVX1 U10375 ( .A(n13516), .Y(n13525) );
  NAND3X1 U10376 ( .A(\forney/m1/added [3]), .B(n13513), .C(n10649), .Y(n13495) );
  NOR2X1 U10377 ( .A(\forney/m1/added [1]), .B(n13495), .Y(n13503) );
  NAND3X1 U10378 ( .A(n13504), .B(n13513), .C(n10649), .Y(n13511) );
  INVX1 U10379 ( .A(\forney/m1/added [2]), .Y(n13507) );
  OAI21X1 U10380 ( .A(\add_x_20/n1 ), .B(\forney/m1/added [4]), .C(
        \forney/m1/added [3]), .Y(n13497) );
  NAND2X1 U10381 ( .A(n13507), .B(n13497), .Y(n13519) );
  NAND2X1 U10382 ( .A(n11197), .B(n13504), .Y(n13498) );
  NAND2X1 U10383 ( .A(\forney/m1/added [2]), .B(n13498), .Y(n13502) );
  NAND2X1 U10384 ( .A(n13519), .B(n13502), .Y(n13499) );
  INVX1 U10385 ( .A(\forney/m1/added [1]), .Y(n13506) );
  AOI21X1 U10386 ( .A(n10459), .B(n13499), .C(n13506), .Y(n13520) );
  OR2X1 U10387 ( .A(n13503), .B(n13520), .Y(n13500) );
  AOI21X1 U10388 ( .A(\forney/m1/added [2]), .B(n13525), .C(n13500), .Y(n13533) );
  NAND3X1 U10389 ( .A(\forney/m1/added [3]), .B(\forney/m1/added [4]), .C(
        \add_x_20/n1 ), .Y(n13508) );
  OAI21X1 U10390 ( .A(n13503), .B(n13502), .C(n10872), .Y(n13523) );
  NAND2X1 U10391 ( .A(\forney/m1/added [1]), .B(\forney/m1/added [2]), .Y(
        n13518) );
  INVX1 U10392 ( .A(n13518), .Y(n13505) );
  AOI22X1 U10393 ( .A(n13505), .B(n10615), .C(n11197), .D(n13504), .Y(n13509)
         );
  NAND2X1 U10394 ( .A(n13506), .B(n10459), .Y(n13527) );
  NAND2X1 U10395 ( .A(n13509), .B(n13527), .Y(n13521) );
  NAND2X1 U10396 ( .A(n13523), .B(n13521), .Y(n13531) );
  OR2X1 U10397 ( .A(n10615), .B(n13507), .Y(n13514) );
  OAI21X1 U10398 ( .A(\forney/m1/added [1]), .B(n13514), .C(n13509), .Y(n13510) );
  INVX1 U10399 ( .A(n13510), .Y(n13522) );
  OR2X1 U10400 ( .A(n13531), .B(n13522), .Y(n13552) );
  INVX1 U10401 ( .A(n10459), .Y(n13512) );
  AOI22X1 U10402 ( .A(\forney/m1/added [1]), .B(n11197), .C(n13512), .D(
        \forney/m1/added [2]), .Y(n13515) );
  NAND3X1 U10403 ( .A(n13516), .B(n13515), .C(n13514), .Y(n13517) );
  HAX1 U10404 ( .A(n13552), .B(n13542), .YS(n13528) );
  INVX1 U10405 ( .A(n13521), .Y(n13526) );
  NAND2X1 U10406 ( .A(n13523), .B(n13522), .Y(n13524) );
  AOI21X1 U10407 ( .A(n13526), .B(n13525), .C(n13524), .Y(n13543) );
  OAI21X1 U10408 ( .A(n10540), .B(n13528), .C(n11108), .Y(n13536) );
  HAX1 U10409 ( .A(n13536), .B(n10655), .YS(n13659) );
  INVX1 U10410 ( .A(n10456), .Y(n13545) );
  INVX1 U10411 ( .A(n13542), .Y(n13532) );
  OAI21X1 U10412 ( .A(n11140), .B(n10782), .C(n13532), .Y(n13534) );
  INVX1 U10413 ( .A(n10540), .Y(n13555) );
  AOI22X1 U10414 ( .A(n10782), .B(n11140), .C(n13534), .D(n10429), .Y(n13564)
         );
  NAND2X1 U10415 ( .A(n13536), .B(n13535), .Y(n13537) );
  NOR2X1 U10416 ( .A(n13537), .B(n11162), .Y(n13561) );
  NAND2X1 U10417 ( .A(n11162), .B(n13537), .Y(n13562) );
  OAI21X1 U10418 ( .A(n10525), .B(n13561), .C(n13562), .Y(n13544) );
  OR2X1 U10419 ( .A(n13545), .B(n13544), .Y(n13557) );
  INVX1 U10420 ( .A(n13557), .Y(n13546) );
  AOI22X1 U10421 ( .A(n10624), .B(n13542), .C(n10429), .D(n13540), .Y(n13560)
         );
  OAI21X1 U10422 ( .A(n13546), .B(n10648), .C(n11017), .Y(n13550) );
  AOI21X1 U10423 ( .A(n13550), .B(n13549), .C(n11158), .Y(n13567) );
  OAI21X1 U10424 ( .A(n13550), .B(n13549), .C(n13547), .Y(n13548) );
  AOI21X1 U10425 ( .A(n13550), .B(n13549), .C(n13548), .Y(n13566) );
  NAND2X1 U10426 ( .A(n13552), .B(n11108), .Y(n13554) );
  AOI21X1 U10427 ( .A(n13555), .B(n13554), .C(n10782), .Y(n13569) );
  NAND2X1 U10428 ( .A(n10531), .B(n10647), .Y(n13556) );
  NAND3X1 U10429 ( .A(n13547), .B(n11017), .C(n13557), .Y(n13559) );
  HAX1 U10430 ( .A(n10648), .B(n13559), .YS(n13618) );
  INVX1 U10431 ( .A(n13618), .Y(n13637) );
  INVX1 U10432 ( .A(n13561), .Y(n13563) );
  NAND3X1 U10433 ( .A(n13547), .B(n13563), .C(n13562), .Y(n13565) );
  HAX1 U10434 ( .A(n13565), .B(n10525), .YS(n13640) );
  HAX1 U10435 ( .A(n10531), .B(n10647), .YS(n13615) );
  OAI21X1 U10436 ( .A(n13643), .B(n13637), .C(n11097), .Y(n13657) );
  INVX1 U10437 ( .A(n13640), .Y(n13619) );
  INVX1 U10438 ( .A(n13567), .Y(n13568) );
  OAI21X1 U10439 ( .A(n13638), .B(n13618), .C(n13643), .Y(n13570) );
  NAND3X1 U10440 ( .A(n13571), .B(n13570), .C(n13659), .Y(n13572) );
  OAI21X1 U10441 ( .A(n13659), .B(n13657), .C(n13572), .Y(n13573) );
  INVX1 U10442 ( .A(n13574), .Y(n13754) );
  NAND3X1 U10443 ( .A(n13575), .B(n10609), .C(n10742), .Y(n13578) );
  INVX1 U10444 ( .A(n13576), .Y(n13577) );
  AOI22X1 U10445 ( .A(n13888), .B(n13578), .C(n13694), .D(n13577), .Y(n13583)
         );
  AOI21X1 U10446 ( .A(n13580), .B(n13684), .C(n13579), .Y(n13581) );
  OAI21X1 U10447 ( .A(n13583), .B(n11172), .C(n13581), .Y(n13584) );
  OAI21X1 U10448 ( .A(n13695), .B(n13754), .C(n13584), .Y(n13748) );
  NAND2X1 U10449 ( .A(n13586), .B(n10609), .Y(n13587) );
  AOI22X1 U10450 ( .A(n12827), .B(n13589), .C(n11203), .D(n13587), .Y(n13890)
         );
  NAND2X1 U10451 ( .A(n13591), .B(n10798), .Y(n13892) );
  NAND3X1 U10452 ( .A(n13890), .B(n11195), .C(n13892), .Y(n13595) );
  MUX2X1 U10453 ( .B(n11210), .A(n13592), .S(n13489), .Y(n13594) );
  AOI22X1 U10454 ( .A(n13752), .B(n13595), .C(n13594), .D(n10664), .Y(n13597)
         );
  NAND2X1 U10455 ( .A(n13597), .B(n13596), .Y(n13598) );
  AOI21X1 U10456 ( .A(n10698), .B(n13753), .C(n13599), .Y(n13749) );
  INVX1 U10457 ( .A(n11175), .Y(n13675) );
  OAI21X1 U10458 ( .A(n13602), .B(n13752), .C(n13601), .Y(n13745) );
  AOI22X1 U10459 ( .A(n11228), .B(n10632), .C(n10636), .D(n13745), .Y(n13603)
         );
  MUX2X1 U10460 ( .B(msg[43]), .A(n13604), .S(n13603), .Y(decoded[43]) );
  INVX1 U10461 ( .A(n13627), .Y(n13606) );
  NAND2X1 U10462 ( .A(n13606), .B(n13628), .Y(n13608) );
  AOI22X1 U10463 ( .A(n13605), .B(n13608), .C(n13606), .D(n13626), .Y(n13611)
         );
  OAI21X1 U10464 ( .A(n13631), .B(n10418), .C(n13607), .Y(n13612) );
  INVX1 U10465 ( .A(n13608), .Y(n13610) );
  AOI22X1 U10466 ( .A(n13610), .B(n13626), .C(n13627), .D(n13609), .Y(n13649)
         );
  AOI22X1 U10467 ( .A(n10863), .B(n11142), .C(n10418), .D(n13631), .Y(n13633)
         );
  INVX1 U10468 ( .A(n11208), .Y(n13648) );
  AOI22X1 U10469 ( .A(n11208), .B(n13612), .C(n10395), .D(n13648), .Y(n13613)
         );
  NOR2X1 U10470 ( .A(n13640), .B(n13637), .Y(n13614) );
  INVX1 U10471 ( .A(n13615), .Y(n13636) );
  AOI22X1 U10472 ( .A(n13615), .B(n13614), .C(n13637), .D(n13636), .Y(n13621)
         );
  NOR2X1 U10473 ( .A(n13659), .B(n13638), .Y(n13616) );
  AOI22X1 U10474 ( .A(n10410), .B(n13659), .C(n13618), .D(n13616), .Y(n13622)
         );
  NAND3X1 U10475 ( .A(n13636), .B(n13619), .C(n13618), .Y(n13617) );
  OAI21X1 U10476 ( .A(n13619), .B(n13618), .C(n13617), .Y(n13658) );
  INVX1 U10477 ( .A(n13659), .Y(n13620) );
  AOI22X1 U10478 ( .A(n13659), .B(n13658), .C(n10410), .D(n13620), .Y(n13642)
         );
  AOI22X1 U10479 ( .A(n13643), .B(n13622), .C(n10419), .D(n10633), .Y(n13623)
         );
  AOI22X1 U10480 ( .A(n10711), .B(n11228), .C(n10704), .D(n13745), .Y(n13624)
         );
  MUX2X1 U10481 ( .B(msg[42]), .A(n13625), .S(n13624), .Y(decoded[42]) );
  NAND3X1 U10482 ( .A(n13628), .B(n13627), .C(n13626), .Y(n13629) );
  NAND3X1 U10483 ( .A(n13648), .B(n10811), .C(n13629), .Y(n13647) );
  AOI22X1 U10484 ( .A(n10863), .B(n13647), .C(n11142), .D(n13631), .Y(n13632)
         );
  AOI21X1 U10485 ( .A(n11208), .B(n10395), .C(n13632), .Y(n13635) );
  NAND2X1 U10486 ( .A(n13637), .B(n13636), .Y(n13639) );
  OAI21X1 U10487 ( .A(n13640), .B(n13639), .C(n11097), .Y(n13655) );
  AOI21X1 U10488 ( .A(n13659), .B(n13655), .C(n13643), .Y(n13656) );
  OAI21X1 U10489 ( .A(n13659), .B(n13658), .C(n13656), .Y(n13641) );
  OAI21X1 U10490 ( .A(n10633), .B(n10419), .C(n13641), .Y(n13644) );
  AOI22X1 U10491 ( .A(n10712), .B(n11228), .C(n10705), .D(n13745), .Y(n13645)
         );
  MUX2X1 U10492 ( .B(msg[41]), .A(n13646), .S(n13645), .Y(decoded[41]) );
  OAI21X1 U10493 ( .A(n11142), .B(n13648), .C(n13647), .Y(n13653) );
  AOI21X1 U10494 ( .A(n13651), .B(n10863), .C(n13650), .Y(n13652) );
  OAI21X1 U10495 ( .A(n10863), .B(n13653), .C(n13652), .Y(n13713) );
  AOI22X1 U10496 ( .A(n13659), .B(n13657), .C(n13656), .D(n13655), .Y(n13663)
         );
  NOR2X1 U10497 ( .A(n13659), .B(n13658), .Y(n13660) );
  AOI22X1 U10498 ( .A(n10713), .B(n11228), .C(n10706), .D(n13745), .Y(n13665)
         );
  MUX2X1 U10499 ( .B(msg[40]), .A(n13666), .S(n13665), .Y(decoded[40]) );
  NOR3X1 U10500 ( .A(n10728), .B(n13748), .C(n13675), .Y(n13789) );
  AOI22X1 U10501 ( .A(n10714), .B(n11228), .C(n13789), .D(n13745), .Y(n13668)
         );
  MUX2X1 U10502 ( .B(msg[39]), .A(n13669), .S(n13668), .Y(decoded[39]) );
  NOR3X1 U10503 ( .A(n13748), .B(n13675), .C(n11170), .Y(n13793) );
  AOI22X1 U10504 ( .A(n10715), .B(n11228), .C(n13793), .D(n13745), .Y(n13670)
         );
  MUX2X1 U10505 ( .B(msg[38]), .A(n13671), .S(n13670), .Y(decoded[38]) );
  NOR3X1 U10506 ( .A(n13748), .B(n13675), .C(n10740), .Y(n13797) );
  AOI22X1 U10507 ( .A(n10716), .B(n11228), .C(n13797), .D(n13745), .Y(n13672)
         );
  MUX2X1 U10508 ( .B(msg[37]), .A(n13673), .S(n13672), .Y(decoded[37]) );
  NOR3X1 U10509 ( .A(n13748), .B(n13675), .C(n13712), .Y(n13801) );
  AOI22X1 U10510 ( .A(n10717), .B(n11228), .C(n13801), .D(n13745), .Y(n13676)
         );
  MUX2X1 U10511 ( .B(msg[36]), .A(n13677), .S(n13676), .Y(decoded[36]) );
  NOR3X1 U10512 ( .A(n13684), .B(n13753), .C(n13702), .Y(n13804) );
  AOI22X1 U10513 ( .A(n13804), .B(n11228), .C(n10707), .D(n13745), .Y(n13678)
         );
  MUX2X1 U10514 ( .B(msg[35]), .A(n13679), .S(n13678), .Y(decoded[35]) );
  NOR3X1 U10515 ( .A(n13684), .B(n13753), .C(n13759), .Y(n13808) );
  AOI22X1 U10516 ( .A(n13808), .B(n11228), .C(n10708), .D(n13745), .Y(n13680)
         );
  MUX2X1 U10517 ( .B(msg[34]), .A(n13681), .S(n13680), .Y(decoded[34]) );
  NOR3X1 U10518 ( .A(n13684), .B(n13753), .C(n13762), .Y(n13812) );
  AOI22X1 U10519 ( .A(n13812), .B(n11228), .C(n10709), .D(n13745), .Y(n13682)
         );
  MUX2X1 U10520 ( .B(msg[33]), .A(n13683), .S(n13682), .Y(decoded[33]) );
  NOR3X1 U10521 ( .A(n13684), .B(n13753), .C(n13713), .Y(n13817) );
  AOI22X1 U10522 ( .A(n13817), .B(n11228), .C(n10710), .D(n13745), .Y(n13687)
         );
  MUX2X1 U10523 ( .B(msg[32]), .A(n13688), .S(n13687), .Y(decoded[32]) );
  NAND3X1 U10524 ( .A(n13692), .B(n11195), .C(n10742), .Y(n13701) );
  AOI22X1 U10525 ( .A(n13752), .B(n11198), .C(n13694), .D(n13693), .Y(n13699)
         );
  NAND2X1 U10526 ( .A(n13697), .B(n10477), .Y(n13906) );
  INVX1 U10527 ( .A(n13906), .Y(n13898) );
  NAND3X1 U10528 ( .A(n13903), .B(n13898), .C(n13888), .Y(n13698) );
  NAND2X1 U10529 ( .A(n13699), .B(n13698), .Y(n13700) );
  AOI22X1 U10530 ( .A(n13752), .B(n13701), .C(n10665), .D(n13700), .Y(n13747)
         );
  NOR3X1 U10531 ( .A(n11175), .B(n13748), .C(n13741), .Y(n13715) );
  INVX1 U10532 ( .A(n13702), .Y(n13756) );
  NOR3X1 U10533 ( .A(n13750), .B(n13751), .C(n10833), .Y(n13740) );
  NAND3X1 U10534 ( .A(n13754), .B(n13753), .C(n13740), .Y(n13703) );
  INVX1 U10535 ( .A(n13703), .Y(n13714) );
  AOI22X1 U10536 ( .A(n13689), .B(n13715), .C(n13756), .D(n13714), .Y(n13704)
         );
  MUX2X1 U10537 ( .B(msg[31]), .A(n13705), .S(n13704), .Y(decoded[31]) );
  AOI22X1 U10538 ( .A(n13706), .B(n13715), .C(n10638), .D(n13714), .Y(n13707)
         );
  MUX2X1 U10539 ( .B(msg[30]), .A(n13708), .S(n13707), .Y(decoded[30]) );
  AOI22X1 U10540 ( .A(n13709), .B(n13715), .C(n10639), .D(n13714), .Y(n13710)
         );
  MUX2X1 U10541 ( .B(msg[29]), .A(n13711), .S(n13710), .Y(decoded[29]) );
  INVX1 U10542 ( .A(n13712), .Y(n13768) );
  INVX1 U10543 ( .A(n13713), .Y(n13766) );
  AOI22X1 U10544 ( .A(n13768), .B(n13715), .C(n13766), .D(n13714), .Y(n13716)
         );
  MUX2X1 U10545 ( .B(msg[28]), .A(n13717), .S(n13716), .Y(decoded[28]) );
  AOI22X1 U10546 ( .A(n10636), .B(n11229), .C(n10632), .D(n13740), .Y(n13718)
         );
  MUX2X1 U10547 ( .B(msg[27]), .A(n13719), .S(n13718), .Y(decoded[27]) );
  AOI22X1 U10548 ( .A(n10704), .B(n11229), .C(n10711), .D(n13740), .Y(n13720)
         );
  MUX2X1 U10549 ( .B(msg[26]), .A(n13721), .S(n13720), .Y(decoded[26]) );
  AOI22X1 U10550 ( .A(n10705), .B(n11229), .C(n10712), .D(n13740), .Y(n13722)
         );
  MUX2X1 U10551 ( .B(msg[25]), .A(n13723), .S(n13722), .Y(decoded[25]) );
  AOI22X1 U10552 ( .A(n10706), .B(n11229), .C(n10713), .D(n13740), .Y(n13724)
         );
  MUX2X1 U10553 ( .B(msg[24]), .A(n13725), .S(n13724), .Y(decoded[24]) );
  AOI22X1 U10554 ( .A(n13789), .B(n11229), .C(n10714), .D(n13740), .Y(n13726)
         );
  MUX2X1 U10555 ( .B(msg[23]), .A(n13727), .S(n13726), .Y(decoded[23]) );
  AOI22X1 U10556 ( .A(n13793), .B(n11229), .C(n10715), .D(n13740), .Y(n13728)
         );
  MUX2X1 U10557 ( .B(msg[22]), .A(n13729), .S(n13728), .Y(decoded[22]) );
  AOI22X1 U10558 ( .A(n13797), .B(n11229), .C(n10716), .D(n13740), .Y(n13730)
         );
  MUX2X1 U10559 ( .B(msg[21]), .A(n13731), .S(n13730), .Y(decoded[21]) );
  AOI22X1 U10560 ( .A(n13801), .B(n11229), .C(n10717), .D(n13740), .Y(n13732)
         );
  MUX2X1 U10561 ( .B(msg[20]), .A(n13733), .S(n13732), .Y(decoded[20]) );
  AOI22X1 U10562 ( .A(n10707), .B(n11229), .C(n13804), .D(n13740), .Y(n13734)
         );
  MUX2X1 U10563 ( .B(msg[19]), .A(n13735), .S(n13734), .Y(decoded[19]) );
  AOI22X1 U10564 ( .A(n10708), .B(n11229), .C(n13808), .D(n13740), .Y(n13736)
         );
  MUX2X1 U10565 ( .B(msg[18]), .A(n13737), .S(n13736), .Y(decoded[18]) );
  AOI22X1 U10566 ( .A(n10709), .B(n11229), .C(n13812), .D(n13740), .Y(n13738)
         );
  MUX2X1 U10567 ( .B(msg[17]), .A(n13739), .S(n13738), .Y(decoded[17]) );
  AOI22X1 U10568 ( .A(n10710), .B(n11229), .C(n13817), .D(n13740), .Y(n13742)
         );
  MUX2X1 U10569 ( .B(msg[16]), .A(n13743), .S(n13742), .Y(decoded[16]) );
  NOR2X1 U10570 ( .A(n13745), .B(n10753), .Y(n13746) );
  NAND2X1 U10571 ( .A(n13747), .B(n13746), .Y(n13771) );
  NOR3X1 U10572 ( .A(n11175), .B(n13748), .C(n13771), .Y(n13767) );
  NOR3X1 U10573 ( .A(n10833), .B(n13751), .C(n10665), .Y(n13816) );
  NAND3X1 U10574 ( .A(n13754), .B(n13753), .C(n13816), .Y(n13755) );
  INVX1 U10575 ( .A(n13755), .Y(n13765) );
  AOI22X1 U10576 ( .A(n13689), .B(n13767), .C(n13756), .D(n13765), .Y(n13757)
         );
  MUX2X1 U10577 ( .B(msg[15]), .A(n13758), .S(n13757), .Y(decoded[15]) );
  AOI22X1 U10578 ( .A(n13706), .B(n13767), .C(n10638), .D(n13765), .Y(n13760)
         );
  MUX2X1 U10579 ( .B(msg[14]), .A(n13761), .S(n13760), .Y(decoded[14]) );
  AOI22X1 U10580 ( .A(n13709), .B(n13767), .C(n10639), .D(n13765), .Y(n13763)
         );
  MUX2X1 U10581 ( .B(msg[13]), .A(n13764), .S(n13763), .Y(decoded[13]) );
  AOI22X1 U10582 ( .A(n13768), .B(n13767), .C(n13766), .D(n13765), .Y(n13769)
         );
  MUX2X1 U10583 ( .B(msg[12]), .A(n13770), .S(n13769), .Y(decoded[12]) );
  INVX1 U10584 ( .A(n13771), .Y(n13818) );
  MUX2X1 U10585 ( .B(msg[11]), .A(n13775), .S(n10974), .Y(decoded[11]) );
  AOI22X1 U10586 ( .A(n10704), .B(n13818), .C(n10711), .D(n13816), .Y(n13778)
         );
  MUX2X1 U10587 ( .B(msg[10]), .A(n13779), .S(n13778), .Y(decoded[10]) );
  AOI22X1 U10588 ( .A(n10705), .B(n13818), .C(n10712), .D(n13816), .Y(n13782)
         );
  MUX2X1 U10589 ( .B(msg[9]), .A(n13783), .S(n13782), .Y(decoded[9]) );
  AOI22X1 U10590 ( .A(n10706), .B(n13818), .C(n10713), .D(n13816), .Y(n13786)
         );
  MUX2X1 U10591 ( .B(msg[8]), .A(n13787), .S(n13786), .Y(decoded[8]) );
  AOI22X1 U10592 ( .A(n13789), .B(n13818), .C(n10714), .D(n13816), .Y(n13790)
         );
  MUX2X1 U10593 ( .B(msg[7]), .A(n13791), .S(n13790), .Y(decoded[7]) );
  AOI22X1 U10594 ( .A(n13793), .B(n13818), .C(n10715), .D(n13816), .Y(n13794)
         );
  MUX2X1 U10595 ( .B(msg[6]), .A(n13795), .S(n13794), .Y(decoded[6]) );
  AOI22X1 U10596 ( .A(n13797), .B(n13818), .C(n10716), .D(n13816), .Y(n13798)
         );
  MUX2X1 U10597 ( .B(msg[5]), .A(n13799), .S(n13798), .Y(decoded[5]) );
  AOI22X1 U10598 ( .A(n13801), .B(n13818), .C(n10717), .D(n13816), .Y(n13802)
         );
  MUX2X1 U10599 ( .B(msg[4]), .A(n13803), .S(n13802), .Y(decoded[4]) );
  AOI22X1 U10600 ( .A(n10707), .B(n13818), .C(n13804), .D(n13816), .Y(n13806)
         );
  MUX2X1 U10601 ( .B(msg[3]), .A(n13807), .S(n13806), .Y(decoded[3]) );
  AOI22X1 U10602 ( .A(n10708), .B(n13818), .C(n13808), .D(n13816), .Y(n13810)
         );
  MUX2X1 U10603 ( .B(msg[2]), .A(n13811), .S(n13810), .Y(decoded[2]) );
  AOI22X1 U10604 ( .A(n10709), .B(n13818), .C(n13812), .D(n13816), .Y(n13814)
         );
  MUX2X1 U10605 ( .B(msg[1]), .A(n13815), .S(n13814), .Y(decoded[1]) );
  AOI22X1 U10606 ( .A(n10710), .B(n13818), .C(n13817), .D(n13816), .Y(n13820)
         );
  MUX2X1 U10607 ( .B(msg[0]), .A(n13821), .S(n13820), .Y(decoded[0]) );
  AND2X1 U10608 ( .A(n13823), .B(n10501), .Y(n13825) );
  OAI21X1 U10609 ( .A(n13826), .B(n13825), .C(n11127), .Y(n10380) );
  OAI21X1 U10610 ( .A(n13830), .B(n13829), .C(n11137), .Y(n10374) );
  NAND2X1 U10611 ( .A(n13831), .B(n13830), .Y(n13832) );
  MUX2X1 U10612 ( .B(n13834), .A(n11137), .S(n13832), .Y(n13835) );
  AOI21X1 U10613 ( .A(n13837), .B(n13836), .C(n13835), .Y(n10373) );
  AOI21X1 U10614 ( .A(n13850), .B(n13852), .C(n10489), .Y(n13839) );
  NAND2X1 U10615 ( .A(n13850), .B(n13854), .Y(n13847) );
  AOI21X1 U10616 ( .A(n13858), .B(n13857), .C(n13847), .Y(n13838) );
  NOR3X1 U10617 ( .A(n13840), .B(n13839), .C(n10967), .Y(
        \lamb/scale_bs2/genblk1[1].mult/added[3] ) );
  NAND2X1 U10618 ( .A(n13842), .B(n13841), .Y(n13843) );
  OAI21X1 U10619 ( .A(n13845), .B(n13844), .C(n13843), .Y(n10370) );
  NAND2X1 U10620 ( .A(n13846), .B(n13848), .Y(n13856) );
  OAI21X1 U10621 ( .A(n13862), .B(n13852), .C(n10489), .Y(
        \lamb/scale_bs2/genblk1[1].mult/added[1] ) );
  OAI21X1 U10622 ( .A(n13848), .B(n13852), .C(n13858), .Y(n13853) );
  NAND2X1 U10623 ( .A(n13850), .B(n10489), .Y(n13851) );
  AOI22X1 U10624 ( .A(n13854), .B(n13853), .C(n13852), .D(n13851), .Y(
        \lamb/scale_bs2/genblk1[1].mult/added[2] ) );
  NAND2X1 U10625 ( .A(n13857), .B(n13855), .Y(n13861) );
  INVX1 U10626 ( .A(n13856), .Y(n13860) );
  NAND2X1 U10627 ( .A(n13858), .B(n13857), .Y(n13859) );
  AOI22X1 U10628 ( .A(n13862), .B(n13861), .C(n13860), .D(n13859), .Y(
        \lamb/scale_bs2/genblk1[1].mult/added[4] ) );
  NAND2X1 U10629 ( .A(n13864), .B(n13863), .Y(n13865) );
  AOI21X1 U10630 ( .A(n13867), .B(n11138), .C(n13865), .Y(n10369) );
  NAND3X1 U10631 ( .A(n10816), .B(n10732), .C(n13868), .Y(n13870) );
  OAI21X1 U10632 ( .A(n13875), .B(n13874), .C(n10626), .Y(n10367) );
  NOR2X1 U10633 ( .A(n13877), .B(n13876), .Y(n13886) );
  AOI21X1 U10634 ( .A(n13880), .B(n13879), .C(n11121), .Y(n13881) );
  INVX1 U10635 ( .A(n13881), .Y(n13883) );
  NAND2X1 U10636 ( .A(n13883), .B(n11054), .Y(n13884) );
  AOI21X1 U10637 ( .A(n13886), .B(n13885), .C(n13884), .Y(n10366) );
  INVX1 U10638 ( .A(n10480), .Y(n13904) );
  AOI22X1 U10639 ( .A(n13888), .B(n13890), .C(n13889), .D(n11210), .Y(n13895)
         );
  NOR2X1 U10640 ( .A(n13892), .B(n13891), .Y(n13894) );
  OAI21X1 U10641 ( .A(n13895), .B(n13894), .C(n13893), .Y(n13900) );
  NAND3X1 U10642 ( .A(n13898), .B(n13897), .C(n13896), .Y(n13899) );
  NAND3X1 U10643 ( .A(n13901), .B(n13900), .C(n13899), .Y(n13902) );
  OAI21X1 U10644 ( .A(n13904), .B(n13903), .C(n13902), .Y(n13911) );
  AOI21X1 U10645 ( .A(n10384), .B(n13906), .C(n13905), .Y(n13909) );
  OAI21X1 U10646 ( .A(n13909), .B(n13908), .C(n10791), .Y(n13910) );
  NAND2X1 U10647 ( .A(n13914), .B(n10646), .Y(n13916) );
  AOI21X1 U10648 ( .A(n13917), .B(n13916), .C(n13915), .Y(n13919) );
  NAND3X1 U10649 ( .A(n13218), .B(n13919), .C(n13918), .Y(n13920) );
  OAI21X1 U10650 ( .A(n13922), .B(n13921), .C(n13920), .Y(n10363) );
  AOI21X1 U10651 ( .A(n13925), .B(n13924), .C(n10468), .Y(n13926) );
  INVX1 U10652 ( .A(n13926), .Y(n13931) );
  OAI21X1 U10653 ( .A(n10745), .B(n10600), .C(n13928), .Y(n13930) );
  OAI21X1 U10654 ( .A(n13932), .B(n13931), .C(n13930), .Y(n10362) );
  OAI21X1 U10655 ( .A(n13935), .B(n13934), .C(n13933), .Y(n13936) );
  NAND2X1 U10656 ( .A(n13937), .B(n13936), .Y(n13938) );
  AOI22X1 U10657 ( .A(n11139), .B(n10407), .C(n10403), .D(n13938), .Y(n10361)
         );
  AND2X1 U10658 ( .A(n13943), .B(n10495), .Y(n13945) );
  OAI21X1 U10659 ( .A(n10832), .B(n13945), .C(n13944), .Y(n10360) );
endmodule


