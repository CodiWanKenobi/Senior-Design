module tb_System_FromFile();

    reg [0:43] in_data;
    reg [0:59] error_mask;
    reg [0:59] modified_data;
    wire [0:43] out_data;
    wire valid;
    
    RS_Top top(in_data, error_mask, out_data, valid);
    
    integer outFile,inFile;

    initial begin
        outFile = $fopen("Output_Data.txt", "w"); //open file for outputting results to
        inFile = $fopen("RS_Input.txt", "r");
        
        while (! $feof(inFile)) begin           //run until reaching end of file
            $fscanf(inFile, "%h", in_data);  //read in a line of the text file
            $fscanf(inFile, "%h", error_mask);  //read in a line of the text file
//            $ferror(inFile,str);
//            $display("%s",str);
            #50
            $fdisplay(outFile, "Input data: %h", in_data);   //write data 
            $fdisplay(outFile, "Error mask: %h", error_mask);   //write data 
            $fdisplay(outFile, "Corrected data: %h", out_data);   //write data 
            if (((in_data == out_data) && valid) || ((in_data != out_data) && (~valid))) begin
                $fdisplay(outFile, "Success\n");   //write data 
            end else begin
                $fdisplay(outFile, "Failure\n");   //write data 
            end
            $fflush(outFile);
            #50;
        end
    end
endmodule

module RS_Top (in, mask, out, valid);
   input  [0:43] in;
   input  [0:59] mask;
   output [0:43] out;
   output valid;
   
   wire [0:59] encoded;
   wire [0:59] masked;
   assign masked = encoded ^ mask;
   RS_Encoder_Optimized enc(in, encoded);
   RS_Decoder dec(masked, out, valid);
endmodule

module RS_Encoder_Optimized ( in, out );
  input [0:43] in;
  output [0:59] out;
  wire   n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439;
  assign out[0] = in[0];
  assign out[1] = in[1];
  assign out[2] = in[2];
  assign out[3] = in[3];
  assign out[4] = in[4];
  assign out[5] = in[5];
  assign out[6] = in[6];
  assign out[7] = in[7];
  assign out[8] = in[8];
  assign out[9] = in[9];
  assign out[10] = in[10];
  assign out[11] = in[11];
  assign out[12] = in[12];
  assign out[13] = in[13];
  assign out[14] = in[14];
  assign out[15] = in[15];
  assign out[16] = in[16];
  assign out[17] = in[17];
  assign out[18] = in[18];
  assign out[19] = in[19];
  assign out[20] = in[20];
  assign out[21] = in[21];
  assign out[22] = in[22];
  assign out[23] = in[23];
  assign out[24] = in[24];
  assign out[25] = in[25];
  assign out[26] = in[26];
  assign out[27] = in[27];
  assign out[28] = in[28];
  assign out[29] = in[29];
  assign out[30] = in[30];
  assign out[31] = in[31];
  assign out[32] = in[32];
  assign out[33] = in[33];
  assign out[34] = in[34];
  assign out[35] = in[35];
  assign out[36] = in[36];
  assign out[37] = in[37];
  assign out[38] = in[38];
  assign out[39] = in[39];
  assign out[40] = in[40];
  assign out[41] = in[41];
  assign out[42] = in[42];
  assign out[43] = in[43];

  BUFX2 U234 ( .A(n248), .Y(n216) );
  BUFX2 U235 ( .A(n260), .Y(n217) );
  BUFX2 U236 ( .A(n280), .Y(n218) );
  BUFX2 U237 ( .A(n382), .Y(n219) );
  BUFX2 U238 ( .A(n396), .Y(n220) );
  BUFX2 U239 ( .A(n426), .Y(n221) );
  BUFX2 U240 ( .A(n298), .Y(n222) );
  BUFX2 U241 ( .A(n367), .Y(n223) );
  BUFX2 U242 ( .A(n282), .Y(n224) );
  BUFX2 U243 ( .A(n337), .Y(n225) );
  BUFX2 U244 ( .A(n289), .Y(n226) );
  BUFX2 U245 ( .A(n432), .Y(n227) );
  BUFX2 U246 ( .A(n263), .Y(n228) );
  BUFX2 U247 ( .A(n267), .Y(n229) );
  BUFX2 U248 ( .A(n325), .Y(n230) );
  BUFX2 U249 ( .A(n410), .Y(n231) );
  BUFX2 U250 ( .A(n276), .Y(n232) );
  BUFX2 U251 ( .A(n319), .Y(n233) );
  BUFX2 U252 ( .A(n368), .Y(n234) );
  BUFX2 U253 ( .A(n372), .Y(n235) );
  BUFX2 U254 ( .A(n322), .Y(n236) );
  BUFX2 U255 ( .A(n427), .Y(n237) );
  INVX1 U256 ( .A(in[23]), .Y(n268) );
  INVX1 U257 ( .A(in[14]), .Y(n424) );
  MUX2X1 U258 ( .B(n424), .A(in[14]), .S(in[38]), .Y(n413) );
  MUX2X1 U259 ( .B(n268), .A(in[23]), .S(n413), .Y(n311) );
  INVX1 U260 ( .A(n311), .Y(n240) );
  INVX1 U261 ( .A(in[31]), .Y(n407) );
  MUX2X1 U262 ( .B(n407), .A(in[31]), .S(in[11]), .Y(n350) );
  INVX1 U263 ( .A(n350), .Y(n238) );
  INVX1 U264 ( .A(in[0]), .Y(n291) );
  MUX2X1 U265 ( .B(n291), .A(in[0]), .S(in[42]), .Y(n313) );
  MUX2X1 U266 ( .B(n238), .A(n350), .S(n313), .Y(n239) );
  MUX2X1 U267 ( .B(n240), .A(n311), .S(n239), .Y(n385) );
  INVX1 U268 ( .A(in[28]), .Y(n315) );
  INVX1 U269 ( .A(in[27]), .Y(n292) );
  AOI22X1 U270 ( .A(in[27]), .B(in[28]), .C(n315), .D(n292), .Y(n427) );
  INVX1 U271 ( .A(n237), .Y(n428) );
  INVX1 U272 ( .A(in[41]), .Y(n394) );
  INVX1 U273 ( .A(in[19]), .Y(n283) );
  AOI22X1 U274 ( .A(in[19]), .B(in[41]), .C(n394), .D(n283), .Y(n289) );
  MUX2X1 U275 ( .B(n428), .A(n237), .S(n226), .Y(n246) );
  INVX1 U276 ( .A(in[7]), .Y(n383) );
  INVX1 U277 ( .A(in[26]), .Y(n330) );
  INVX1 U278 ( .A(in[5]), .Y(n341) );
  INVX1 U279 ( .A(in[12]), .Y(n374) );
  AOI22X1 U280 ( .A(in[12]), .B(in[5]), .C(n341), .D(n374), .Y(n276) );
  MUX2X1 U281 ( .B(n330), .A(in[26]), .S(n232), .Y(n241) );
  MUX2X1 U282 ( .B(n383), .A(in[7]), .S(n241), .Y(n252) );
  INVX1 U283 ( .A(in[2]), .Y(n284) );
  INVX1 U284 ( .A(in[24]), .Y(n257) );
  INVX1 U285 ( .A(in[20]), .Y(n336) );
  MUX2X1 U286 ( .B(n336), .A(in[20]), .S(in[18]), .Y(n258) );
  MUX2X1 U287 ( .B(n257), .A(in[24]), .S(n258), .Y(n242) );
  MUX2X1 U288 ( .B(n284), .A(in[2]), .S(n242), .Y(n274) );
  INVX1 U289 ( .A(in[33]), .Y(n390) );
  INVX1 U290 ( .A(in[8]), .Y(n338) );
  INVX1 U291 ( .A(in[25]), .Y(n279) );
  INVX1 U292 ( .A(in[17]), .Y(n397) );
  INVX1 U293 ( .A(in[32]), .Y(n278) );
  AOI22X1 U294 ( .A(in[32]), .B(in[17]), .C(n397), .D(n278), .Y(n267) );
  MUX2X1 U295 ( .B(n279), .A(in[25]), .S(n229), .Y(n415) );
  MUX2X1 U296 ( .B(n338), .A(in[8]), .S(n415), .Y(n243) );
  MUX2X1 U297 ( .B(n390), .A(in[33]), .S(n243), .Y(n244) );
  FAX1 U298 ( .A(n252), .B(n274), .C(n244), .YS(n245) );
  FAX1 U299 ( .A(n385), .B(n246), .C(n245), .YS(out[59]) );
  INVX1 U300 ( .A(in[30]), .Y(n430) );
  INVX1 U301 ( .A(in[35]), .Y(n423) );
  AOI22X1 U302 ( .A(in[35]), .B(in[2]), .C(n284), .D(n423), .Y(n298) );
  MUX2X1 U303 ( .B(n430), .A(in[30]), .S(n222), .Y(n256) );
  INVX1 U304 ( .A(n256), .Y(n247) );
  INVX1 U305 ( .A(in[40]), .Y(n302) );
  AOI22X1 U306 ( .A(in[33]), .B(in[40]), .C(n302), .D(n390), .Y(n367) );
  MUX2X1 U307 ( .B(n256), .A(n247), .S(n223), .Y(n310) );
  INVX1 U308 ( .A(n310), .Y(n255) );
  MUX2X1 U309 ( .B(n268), .A(in[23]), .S(n226), .Y(n420) );
  INVX1 U310 ( .A(in[13]), .Y(n293) );
  MUX2X1 U311 ( .B(n293), .A(in[13]), .S(n237), .Y(n362) );
  INVX1 U312 ( .A(in[21]), .Y(n317) );
  INVX1 U313 ( .A(in[16]), .Y(n314) );
  INVX1 U314 ( .A(in[37]), .Y(n290) );
  INVX1 U315 ( .A(in[3]), .Y(n406) );
  AOI22X1 U316 ( .A(in[3]), .B(in[8]), .C(n338), .D(n406), .Y(n368) );
  MUX2X1 U317 ( .B(n290), .A(in[37]), .S(n234), .Y(n353) );
  MUX2X1 U318 ( .B(n314), .A(in[16]), .S(n353), .Y(n405) );
  MUX2X1 U319 ( .B(n317), .A(in[21]), .S(n405), .Y(n288) );
  INVX1 U320 ( .A(in[18]), .Y(n249) );
  INVX1 U321 ( .A(in[36]), .Y(n277) );
  AOI22X1 U322 ( .A(in[36]), .B(in[0]), .C(n291), .D(n277), .Y(n248) );
  MUX2X1 U323 ( .B(n249), .A(in[18]), .S(n216), .Y(n250) );
  MUX2X1 U324 ( .B(n257), .A(in[24]), .S(n250), .Y(n251) );
  FAX1 U325 ( .A(n288), .B(n252), .C(n251), .YS(n253) );
  FAX1 U326 ( .A(n420), .B(n362), .C(n253), .YS(n254) );
  MUX2X1 U327 ( .B(n310), .A(n255), .S(n254), .Y(out[48]) );
  INVX1 U328 ( .A(in[9]), .Y(n266) );
  MUX2X1 U329 ( .B(n266), .A(in[9]), .S(n256), .Y(n294) );
  INVX1 U330 ( .A(in[4]), .Y(n335) );
  AOI22X1 U331 ( .A(in[4]), .B(in[26]), .C(n330), .D(n335), .Y(n282) );
  MUX2X1 U332 ( .B(n383), .A(in[7]), .S(n224), .Y(n392) );
  INVX1 U333 ( .A(n392), .Y(n393) );
  AOI22X1 U334 ( .A(n392), .B(in[24]), .C(n257), .D(n393), .Y(n319) );
  INVX1 U335 ( .A(in[39]), .Y(n421) );
  MUX2X1 U336 ( .B(n421), .A(in[39]), .S(n258), .Y(n381) );
  INVX1 U337 ( .A(n381), .Y(n380) );
  AOI22X1 U338 ( .A(n381), .B(in[25]), .C(n279), .D(n380), .Y(n325) );
  INVX1 U339 ( .A(in[1]), .Y(n408) );
  MUX2X1 U340 ( .B(n408), .A(in[1]), .S(in[43]), .Y(n265) );
  INVX1 U341 ( .A(n265), .Y(n259) );
  MUX2X1 U342 ( .B(n265), .A(n259), .S(n350), .Y(n339) );
  XNOR2X1 U343 ( .A(n230), .B(n339), .Y(n306) );
  INVX1 U344 ( .A(in[15]), .Y(n395) );
  AOI22X1 U345 ( .A(in[13]), .B(in[15]), .C(n395), .D(n293), .Y(n263) );
  INVX1 U346 ( .A(n234), .Y(n369) );
  AOI22X1 U347 ( .A(in[5]), .B(in[36]), .C(n277), .D(n341), .Y(n260) );
  MUX2X1 U348 ( .B(n428), .A(n237), .S(n217), .Y(n261) );
  MUX2X1 U349 ( .B(n369), .A(n234), .S(n261), .Y(n262) );
  FAX1 U350 ( .A(n306), .B(n228), .C(n262), .YS(n264) );
  FAX1 U351 ( .A(n294), .B(n233), .C(n264), .YS(out[55]) );
  INVX1 U352 ( .A(n274), .Y(n275) );
  MUX2X1 U353 ( .B(n317), .A(in[21]), .S(n265), .Y(n365) );
  INVX1 U354 ( .A(n365), .Y(n366) );
  INVX1 U355 ( .A(in[6]), .Y(n351) );
  AOI22X1 U356 ( .A(in[9]), .B(in[6]), .C(n351), .D(n266), .Y(n322) );
  MUX2X1 U357 ( .B(n430), .A(in[30]), .S(n236), .Y(n401) );
  MUX2X1 U358 ( .B(n366), .A(n365), .S(n401), .Y(n272) );
  INVX1 U359 ( .A(n353), .Y(n354) );
  MUX2X1 U360 ( .B(n268), .A(in[23]), .S(n229), .Y(n300) );
  MUX2X1 U361 ( .B(n354), .A(n353), .S(n300), .Y(n271) );
  MUX2X1 U362 ( .B(n315), .A(in[28]), .S(n232), .Y(n269) );
  MUX2X1 U363 ( .B(n291), .A(in[0]), .S(n269), .Y(n270) );
  FAX1 U364 ( .A(n272), .B(n271), .C(n270), .YS(n273) );
  MUX2X1 U365 ( .B(n275), .A(n274), .S(n273), .Y(out[46]) );
  INVX1 U366 ( .A(in[10]), .Y(n425) );
  MUX2X1 U367 ( .B(n425), .A(in[10]), .S(n232), .Y(n348) );
  INVX1 U368 ( .A(in[29]), .Y(n324) );
  AOI22X1 U369 ( .A(in[29]), .B(n277), .C(in[36]), .D(n324), .Y(n372) );
  XNOR2X1 U370 ( .A(n348), .B(n235), .Y(n388) );
  MUX2X1 U371 ( .B(n278), .A(in[32]), .S(n388), .Y(n321) );
  MUX2X1 U372 ( .B(n424), .A(in[14]), .S(n321), .Y(n297) );
  AOI22X1 U373 ( .A(in[25]), .B(in[31]), .C(n407), .D(n279), .Y(n280) );
  MUX2X1 U374 ( .B(n302), .A(in[40]), .S(n218), .Y(n281) );
  MUX2X1 U375 ( .B(n292), .A(in[27]), .S(n281), .Y(n286) );
  MUX2X1 U376 ( .B(n283), .A(in[19]), .S(n224), .Y(n364) );
  MUX2X1 U377 ( .B(n284), .A(in[2]), .S(n364), .Y(n285) );
  FAX1 U378 ( .A(n286), .B(n236), .C(n285), .YS(n287) );
  FAX1 U379 ( .A(n297), .B(n288), .C(n287), .YS(out[52]) );
  INVX1 U380 ( .A(in[34]), .Y(n323) );
  MUX2X1 U381 ( .B(in[34]), .A(n323), .S(n392), .Y(n309) );
  XNOR2X1 U382 ( .A(n365), .B(n309), .Y(n438) );
  MUX2X1 U383 ( .B(n290), .A(in[37]), .S(n226), .Y(n416) );
  MUX2X1 U384 ( .B(n291), .A(in[0]), .S(n416), .Y(n295) );
  INVX1 U385 ( .A(in[22]), .Y(n347) );
  AOI22X1 U386 ( .A(in[27]), .B(in[22]), .C(n347), .D(n292), .Y(n337) );
  MUX2X1 U387 ( .B(n293), .A(in[13]), .S(n225), .Y(n328) );
  FAX1 U388 ( .A(n295), .B(n328), .C(n294), .YS(n296) );
  FAX1 U389 ( .A(n438), .B(n297), .C(n296), .YS(out[57]) );
  INVX1 U390 ( .A(n309), .Y(n308) );
  INVX1 U391 ( .A(n235), .Y(n371) );
  MUX2X1 U392 ( .B(n235), .A(n371), .S(n222), .Y(n345) );
  MUX2X1 U393 ( .B(n351), .A(in[6]), .S(n345), .Y(n299) );
  MUX2X1 U394 ( .B(n374), .A(in[12]), .S(n299), .Y(n305) );
  MUX2X1 U395 ( .B(n395), .A(in[15]), .S(n300), .Y(n301) );
  MUX2X1 U396 ( .B(n302), .A(in[40]), .S(n301), .Y(n303) );
  MUX2X1 U397 ( .B(n347), .A(in[22]), .S(n303), .Y(n304) );
  FAX1 U398 ( .A(n306), .B(n305), .C(n304), .YS(n307) );
  MUX2X1 U399 ( .B(n309), .A(n308), .S(n307), .Y(out[51]) );
  INVX1 U400 ( .A(in[43]), .Y(n312) );
  XNOR2X1 U401 ( .A(n311), .B(n310), .Y(n359) );
  MUX2X1 U402 ( .B(n312), .A(in[43]), .S(n359), .Y(n333) );
  MUX2X1 U403 ( .B(n395), .A(in[15]), .S(n313), .Y(n326) );
  MUX2X1 U404 ( .B(n314), .A(in[16]), .S(n326), .Y(n435) );
  MUX2X1 U405 ( .B(n315), .A(in[28]), .S(n381), .Y(n316) );
  MUX2X1 U406 ( .B(n317), .A(in[21]), .S(n316), .Y(n318) );
  FAX1 U407 ( .A(n435), .B(n233), .C(n318), .YS(n320) );
  FAX1 U408 ( .A(n321), .B(n333), .C(n320), .YS(out[50]) );
  INVX1 U409 ( .A(n333), .Y(n334) );
  MUX2X1 U410 ( .B(n323), .A(in[34]), .S(n236), .Y(n361) );
  MUX2X1 U411 ( .B(n324), .A(in[29]), .S(n361), .Y(n418) );
  INVX1 U412 ( .A(n326), .Y(n327) );
  MUX2X1 U413 ( .B(n327), .A(n326), .S(n230), .Y(n378) );
  MUX2X1 U414 ( .B(n394), .A(in[41]), .S(n328), .Y(n329) );
  MUX2X1 U415 ( .B(n330), .A(in[26]), .S(n329), .Y(n331) );
  FAX1 U416 ( .A(n418), .B(n378), .C(n331), .YS(n332) );
  MUX2X1 U417 ( .B(n334), .A(n333), .S(n332), .Y(out[47]) );
  INVX1 U418 ( .A(n345), .Y(n346) );
  INVX1 U419 ( .A(n435), .Y(n436) );
  AOI22X1 U420 ( .A(in[4]), .B(in[20]), .C(n336), .D(n335), .Y(n410) );
  MUX2X1 U421 ( .B(n436), .A(n435), .S(n231), .Y(n357) );
  MUX2X1 U422 ( .B(n338), .A(in[8]), .S(n225), .Y(n343) );
  MUX2X1 U423 ( .B(in[17]), .A(n397), .S(n339), .Y(n340) );
  MUX2X1 U424 ( .B(n341), .A(in[5]), .S(n340), .Y(n342) );
  FAX1 U425 ( .A(n357), .B(n343), .C(n342), .YS(n344) );
  MUX2X1 U426 ( .B(n346), .A(n345), .S(n344), .Y(out[45]) );
  INVX1 U427 ( .A(n359), .Y(n360) );
  INVX1 U428 ( .A(n348), .Y(n349) );
  MUX2X1 U429 ( .B(n347), .A(in[22]), .S(n362), .Y(n412) );
  MUX2X1 U430 ( .B(n349), .A(n348), .S(n412), .Y(n404) );
  MUX2X1 U431 ( .B(n351), .A(in[6]), .S(n350), .Y(n352) );
  MUX2X1 U432 ( .B(n354), .A(n353), .S(n352), .Y(n355) );
  MUX2X1 U433 ( .B(n408), .A(in[1]), .S(n355), .Y(n356) );
  FAX1 U434 ( .A(n404), .B(n357), .C(n356), .YS(n358) );
  MUX2X1 U435 ( .B(n360), .A(n359), .S(n358), .Y(out[58]) );
  INVX1 U436 ( .A(n378), .Y(n379) );
  INVX1 U437 ( .A(n362), .Y(n363) );
  MUX2X1 U438 ( .B(n363), .A(n362), .S(n361), .Y(n386) );
  MUX2X1 U439 ( .B(n366), .A(n365), .S(n364), .Y(n376) );
  MUX2X1 U440 ( .B(n369), .A(n234), .S(n223), .Y(n370) );
  MUX2X1 U441 ( .B(n235), .A(n371), .S(n370), .Y(n373) );
  MUX2X1 U442 ( .B(n374), .A(in[12]), .S(n373), .Y(n375) );
  FAX1 U443 ( .A(n386), .B(n376), .C(n375), .YS(n377) );
  MUX2X1 U444 ( .B(n379), .A(n378), .S(n377), .Y(out[56]) );
  INVX1 U445 ( .A(n388), .Y(n389) );
  AOI22X1 U446 ( .A(n381), .B(in[17]), .C(n397), .D(n380), .Y(n382) );
  MUX2X1 U447 ( .B(n383), .A(in[7]), .S(n219), .Y(n384) );
  FAX1 U448 ( .A(n386), .B(n385), .C(n384), .YS(n387) );
  MUX2X1 U449 ( .B(n389), .A(n388), .S(n387), .Y(out[54]) );
  MUX2X1 U450 ( .B(n390), .A(in[33]), .S(in[11]), .Y(n391) );
  MUX2X1 U451 ( .B(n393), .A(n392), .S(n391), .Y(n402) );
  INVX1 U452 ( .A(in[38]), .Y(n399) );
  AOI22X1 U453 ( .A(in[41]), .B(in[15]), .C(n395), .D(n394), .Y(n396) );
  MUX2X1 U454 ( .B(n397), .A(in[17]), .S(n220), .Y(n398) );
  MUX2X1 U455 ( .B(n399), .A(in[38]), .S(n398), .Y(n400) );
  FAX1 U456 ( .A(n402), .B(n401), .C(n400), .YS(n403) );
  FAX1 U457 ( .A(n405), .B(n404), .C(n403), .YS(out[53]) );
  INVX1 U458 ( .A(n418), .Y(n419) );
  AOI22X1 U459 ( .A(in[3]), .B(in[31]), .C(n407), .D(n406), .Y(n432) );
  MUX2X1 U460 ( .B(n408), .A(in[1]), .S(in[42]), .Y(n409) );
  FAX1 U461 ( .A(n231), .B(n227), .C(n409), .YS(n411) );
  FAX1 U462 ( .A(n413), .B(n412), .C(n411), .YS(n414) );
  FAX1 U463 ( .A(n416), .B(n415), .C(n414), .YS(n417) );
  MUX2X1 U464 ( .B(n419), .A(n418), .S(n417), .Y(out[49]) );
  INVX1 U465 ( .A(n438), .Y(n439) );
  MUX2X1 U466 ( .B(n421), .A(in[39]), .S(n420), .Y(n422) );
  MUX2X1 U467 ( .B(n423), .A(in[35]), .S(n422), .Y(n433) );
  AOI22X1 U468 ( .A(in[14]), .B(in[10]), .C(n425), .D(n424), .Y(n426) );
  MUX2X1 U469 ( .B(n428), .A(n237), .S(n221), .Y(n429) );
  MUX2X1 U470 ( .B(n430), .A(in[30]), .S(n429), .Y(n431) );
  FAX1 U471 ( .A(n433), .B(n227), .C(n431), .YS(n434) );
  MUX2X1 U472 ( .B(n436), .A(n435), .S(n434), .Y(n437) );
  MUX2X1 U473 ( .B(n439), .A(n438), .S(n437), .Y(out[44]) );
endmodule


module RS_Decoder ( msg, decoded, valid );
  input [0:59] msg;
  output [0:43] decoded;
  output valid;
  wire   \lamb/scale_ts3/genblk1[3].mult/added[1] ,
         \lamb/scale_ts3/genblk1[3].mult/added[2] ,
         \lamb/scale_ts3/genblk1[3].mult/added[3] ,
         \lamb/scale_ts3/genblk1[3].mult/added[4] ,
         \lamb/scale_ts3/genblk1[3].mult/logA[0] ,
         \lamb/scale_ts3/genblk1[3].mult/logA[1] ,
         \lamb/scale_ts3/genblk1[3].mult/logA[2] ,
         \lamb/scale_ts3/genblk1[3].mult/logA[3] ,
         \lamb/scale_ts3/genblk1[2].mult/added[1] ,
         \lamb/scale_ts3/genblk1[2].mult/added[2] ,
         \lamb/scale_ts3/genblk1[2].mult/added[3] ,
         \lamb/scale_ts3/genblk1[2].mult/added[4] ,
         \lamb/scale_ts3/genblk1[2].mult/logA[0] ,
         \lamb/scale_ts3/genblk1[2].mult/logA[1] ,
         \lamb/scale_ts3/genblk1[2].mult/logA[2] ,
         \lamb/scale_ts3/genblk1[2].mult/logA[3] ,
         \lamb/scale_ds3/genblk1[3].mult/added[1] ,
         \lamb/scale_ds3/genblk1[3].mult/added[2] ,
         \lamb/scale_ds3/genblk1[3].mult/added[3] ,
         \lamb/scale_ds3/genblk1[3].mult/added[4] ,
         \lamb/scale_ds3/genblk1[3].mult/logA[0] ,
         \lamb/scale_ds3/genblk1[3].mult/logA[1] ,
         \lamb/scale_ds3/genblk1[3].mult/logA[2] ,
         \lamb/scale_ds3/genblk1[3].mult/logA[3] ,
         \lamb/scale_ds3/genblk1[2].mult/added[1] ,
         \lamb/scale_ds3/genblk1[2].mult/added[2] ,
         \lamb/scale_ds3/genblk1[2].mult/added[3] ,
         \lamb/scale_ds3/genblk1[2].mult/added[4] ,
         \lamb/scale_ds3/genblk1[2].mult/logA[1] ,
         \lamb/scale_ds3/genblk1[2].mult/logA[2] ,
         \lamb/scale_ds3/genblk1[2].mult/logA[3] ,
         \lamb/scale_bs3/genblk1[1].mult/added[1] ,
         \lamb/scale_bs3/genblk1[1].mult/added[2] ,
         \lamb/scale_bs3/genblk1[1].mult/added[3] ,
         \lamb/scale_bs3/genblk1[1].mult/added[4] ,
         \lamb/scale_bs3/genblk1[1].mult/logA[0] ,
         \lamb/scale_bs3/genblk1[1].mult/logA[3] ,
         \lamb/scale_bs3/genblk1[0].mult/added[1] ,
         \lamb/scale_bs3/genblk1[0].mult/added[2] ,
         \lamb/scale_bs3/genblk1[0].mult/added[3] ,
         \lamb/scale_bs3/genblk1[0].mult/added[4] ,
         \lamb/scale_bs3/genblk1[0].mult/logB[0] ,
         \lamb/scale_bs3/genblk1[0].mult/logB[1] ,
         \lamb/scale_bs3/genblk1[0].mult/logB[3] ,
         \lamb/scale_bs3/genblk1[0].mult/logA[0] ,
         \lamb/scale_bs3/genblk1[0].mult/logA[1] ,
         \lamb/scale_bs3/genblk1[0].mult/logA[2] ,
         \lamb/scale_bs3/genblk1[0].mult/logA[3] ,
         \lamb/scale_ls3/genblk1[2].mult/added[1] ,
         \lamb/scale_ls3/genblk1[2].mult/added[2] ,
         \lamb/scale_ls3/genblk1[2].mult/added[3] ,
         \lamb/scale_ls3/genblk1[2].mult/added[4] ,
         \lamb/scale_ls3/genblk1[2].mult/logA[0] ,
         \lamb/scale_ls3/genblk1[2].mult/logA[2] ,
         \lamb/scale_ls3/genblk1[2].mult/logA[3] ,
         \lamb/scale_ls3/genblk1[1].mult/added[1] ,
         \lamb/scale_ls3/genblk1[1].mult/added[2] ,
         \lamb/scale_ls3/genblk1[1].mult/added[3] ,
         \lamb/scale_ls3/genblk1[1].mult/added[4] ,
         \lamb/scale_ls3/genblk1[1].mult/logA[0] ,
         \lamb/scale_ls3/genblk1[1].mult/logA[1] ,
         \lamb/scale_ls3/genblk1[1].mult/logA[2] ,
         \lamb/scale_ls3/genblk1[1].mult/logA[3] ,
         \lamb/scale_ls3/genblk1[0].mult/added[1] ,
         \lamb/scale_ls3/genblk1[0].mult/added[2] ,
         \lamb/scale_ls3/genblk1[0].mult/added[3] ,
         \lamb/scale_ls3/genblk1[0].mult/added[4] ,
         \lamb/scale_ls3/genblk1[0].mult/logB[1] ,
         \lamb/scale_ls3/genblk1[0].mult/logB[2] ,
         \lamb/scale_ls3/genblk1[0].mult/logB[3] ,
         \lamb/scale_ls3/genblk1[0].mult/logA[1] ,
         \lamb/scale_ls3/genblk1[0].mult/logA[2] ,
         \lamb/scale_ls3/genblk1[0].mult/logA[3] ,
         \lamb/scale_ts2/genblk1[3].mult/added[1] ,
         \lamb/scale_ts2/genblk1[3].mult/added[2] ,
         \lamb/scale_ts2/genblk1[3].mult/added[3] ,
         \lamb/scale_ts2/genblk1[3].mult/added[4] ,
         \lamb/scale_ts2/genblk1[3].mult/logA[1] ,
         \lamb/scale_ts2/genblk1[3].mult/logA[2] ,
         \lamb/scale_ts2/genblk1[3].mult/logA[3] ,
         \lamb/scale_ts2/genblk1[2].mult/added[1] ,
         \lamb/scale_ts2/genblk1[2].mult/added[2] ,
         \lamb/scale_ts2/genblk1[2].mult/added[3] ,
         \lamb/scale_ts2/genblk1[2].mult/added[4] ,
         \lamb/scale_ts2/genblk1[2].mult/logA[1] ,
         \lamb/scale_ts2/genblk1[2].mult/logA[2] ,
         \lamb/scale_ts2/genblk1[2].mult/logA[3] ,
         \lamb/scale_ts2/genblk1[1].mult/added[1] ,
         \lamb/scale_ts2/genblk1[1].mult/added[2] ,
         \lamb/scale_ts2/genblk1[1].mult/added[3] ,
         \lamb/scale_ts2/genblk1[1].mult/added[4] ,
         \lamb/scale_ts2/genblk1[1].mult/logA[0] ,
         \lamb/scale_ts2/genblk1[1].mult/logA[1] ,
         \lamb/scale_ts2/genblk1[1].mult/logA[2] ,
         \lamb/scale_ts2/genblk1[1].mult/logA[3] ,
         \lamb/scale_ds2/genblk1[3].mult/added[1] ,
         \lamb/scale_ds2/genblk1[3].mult/added[2] ,
         \lamb/scale_ds2/genblk1[3].mult/added[3] ,
         \lamb/scale_ds2/genblk1[3].mult/added[4] ,
         \lamb/scale_ds2/genblk1[3].mult/logA[0] ,
         \lamb/scale_ds2/genblk1[3].mult/logA[1] ,
         \lamb/scale_ds2/genblk1[3].mult/logA[3] ,
         \lamb/scale_ds2/genblk1[2].mult/added[1] ,
         \lamb/scale_ds2/genblk1[2].mult/added[2] ,
         \lamb/scale_ds2/genblk1[2].mult/added[3] ,
         \lamb/scale_ds2/genblk1[2].mult/added[4] ,
         \lamb/scale_ds2/genblk1[2].mult/logA[0] ,
         \lamb/scale_ds2/genblk1[2].mult/logA[1] ,
         \lamb/scale_ds2/genblk1[2].mult/logA[2] ,
         \lamb/scale_ds2/genblk1[2].mult/logA[3] ,
         \lamb/scale_ds2/genblk1[1].mult/added[1] ,
         \lamb/scale_ds2/genblk1[1].mult/added[2] ,
         \lamb/scale_ds2/genblk1[1].mult/added[3] ,
         \lamb/scale_ds2/genblk1[1].mult/added[4] ,
         \lamb/scale_ds2/genblk1[1].mult/logA[0] ,
         \lamb/scale_ds2/genblk1[1].mult/logA[1] ,
         \lamb/scale_ds2/genblk1[1].mult/logA[2] ,
         \lamb/scale_ds2/genblk1[1].mult/logA[3] ,
         \lamb/scale_bs2/genblk1[1].mult/added[2] ,
         \lamb/scale_bs2/genblk1[1].mult/added[3] ,
         \lamb/scale_bs2/genblk1[1].mult/added[4] ,
         \lamb/scale_bs2/genblk1[0].mult/added[1] ,
         \lamb/scale_bs2/genblk1[0].mult/added[2] ,
         \lamb/scale_bs2/genblk1[0].mult/added[3] ,
         \lamb/scale_bs2/genblk1[0].mult/added[4] ,
         \lamb/scale_bs2/genblk1[0].mult/logA[0] ,
         \lamb/scale_bs2/genblk1[0].mult/logA[2] ,
         \lamb/scale_bs2/genblk1[0].mult/logA[3] ,
         \lamb/scale_ls2/genblk1[2].mult/added[1] ,
         \lamb/scale_ls2/genblk1[2].mult/added[2] ,
         \lamb/scale_ls2/genblk1[2].mult/added[3] ,
         \lamb/scale_ls2/genblk1[2].mult/added[4] ,
         \lamb/scale_ls2/genblk1[1].mult/added[1] ,
         \lamb/scale_ls2/genblk1[1].mult/added[2] ,
         \lamb/scale_ls2/genblk1[1].mult/added[3] ,
         \lamb/scale_ls2/genblk1[1].mult/added[4] ,
         \lamb/scale_ls2/genblk1[1].mult/logA[2] ,
         \lamb/scale_ls2/genblk1[0].mult/added[1] ,
         \lamb/scale_ls2/genblk1[0].mult/added[2] ,
         \lamb/scale_ls2/genblk1[0].mult/added[3] ,
         \lamb/scale_ls2/genblk1[0].mult/added[4] ,
         \lamb/scale_ls2/genblk1[0].mult/logB[0] ,
         \lamb/scale_ls2/genblk1[0].mult/logB[2] ,
         \lamb/scale_ls2/genblk1[0].mult/logA[0] ,
         \lamb/scale_ls2/genblk1[0].mult/logA[1] ,
         \lamb/scale_ls2/genblk1[0].mult/logA[2] ,
         \lamb/scale_ls2/genblk1[0].mult/logA[3] ,
         \lamb/scale_ts1/genblk1[3].mult/added[1] ,
         \lamb/scale_ts1/genblk1[3].mult/added[2] ,
         \lamb/scale_ts1/genblk1[3].mult/added[3] ,
         \lamb/scale_ts1/genblk1[3].mult/added[4] ,
         \lamb/scale_ts1/genblk1[3].mult/logA[0] ,
         \lamb/scale_ts1/genblk1[3].mult/logA[1] ,
         \lamb/scale_ts1/genblk1[2].mult/added[1] ,
         \lamb/scale_ts1/genblk1[2].mult/added[2] ,
         \lamb/scale_ts1/genblk1[2].mult/added[3] ,
         \lamb/scale_ts1/genblk1[2].mult/added[4] ,
         \lamb/scale_ts1/genblk1[2].mult/logA[0] ,
         \lamb/scale_ts1/genblk1[2].mult/logA[1] ,
         \lamb/scale_ts1/genblk1[2].mult/logA[2] ,
         \lamb/scale_ts1/genblk1[1].mult/added[1] ,
         \lamb/scale_ts1/genblk1[1].mult/added[2] ,
         \lamb/scale_ts1/genblk1[1].mult/added[3] ,
         \lamb/scale_ts1/genblk1[1].mult/added[4] ,
         \lamb/scale_ts1/genblk1[1].mult/logA[1] ,
         \lamb/scale_ts1/genblk1[1].mult/logA[3] ,
         \lamb/scale_ts1/genblk1[0].mult/added[1] ,
         \lamb/scale_ts1/genblk1[0].mult/added[2] ,
         \lamb/scale_ts1/genblk1[0].mult/added[3] ,
         \lamb/scale_ts1/genblk1[0].mult/added[4] ,
         \lamb/scale_ts1/genblk1[0].mult/logB[0] ,
         \lamb/scale_ts1/genblk1[0].mult/logB[1] ,
         \lamb/scale_ts1/genblk1[0].mult/logB[2] ,
         \lamb/scale_ts1/genblk1[0].mult/logB[3] ,
         \lamb/scale_ts1/genblk1[0].mult/logA[0] ,
         \lamb/scale_ts1/genblk1[0].mult/logA[1] ,
         \lamb/scale_ts1/genblk1[0].mult/logA[2] ,
         \lamb/scale_ts1/genblk1[0].mult/logA[3] ,
         \lamb/scale_ds1/genblk1[3].mult/added[1] ,
         \lamb/scale_ds1/genblk1[3].mult/added[2] ,
         \lamb/scale_ds1/genblk1[3].mult/added[3] ,
         \lamb/scale_ds1/genblk1[3].mult/added[4] ,
         \lamb/scale_ds1/genblk1[3].mult/logA[2] ,
         \lamb/scale_ds1/genblk1[3].mult/logA[3] ,
         \lamb/scale_ds1/genblk1[2].mult/added[1] ,
         \lamb/scale_ds1/genblk1[2].mult/added[2] ,
         \lamb/scale_ds1/genblk1[2].mult/added[3] ,
         \lamb/scale_ds1/genblk1[2].mult/added[4] ,
         \lamb/scale_ds1/genblk1[2].mult/logA[0] ,
         \lamb/scale_ds1/genblk1[2].mult/logA[3] ,
         \lamb/scale_ds1/genblk1[1].mult/added[1] ,
         \lamb/scale_ds1/genblk1[1].mult/added[2] ,
         \lamb/scale_ds1/genblk1[1].mult/added[3] ,
         \lamb/scale_ds1/genblk1[1].mult/added[4] ,
         \lamb/scale_ds1/genblk1[1].mult/logA[1] ,
         \lamb/scale_ds1/genblk1[1].mult/logA[2] ,
         \lamb/scale_ds1/genblk1[1].mult/logA[3] ,
         \lamb/scale_ls1/genblk1[1].mult/added[2] ,
         \lamb/scale_ls1/genblk1[1].mult/added[3] ,
         \lamb/scale_ts0/genblk1[2].mult/added[1] ,
         \lamb/scale_ts0/genblk1[2].mult/added[2] ,
         \lamb/scale_ts0/genblk1[2].mult/added[3] ,
         \lamb/scale_ts0/genblk1[2].mult/added[4] ,
         \lamb/scale_ts0/genblk1[2].mult/logA[0] ,
         \lamb/scale_ts0/genblk1[2].mult/logA[1] ,
         \lamb/scale_ts0/genblk1[2].mult/logA[3] ,
         \lamb/scale_ts0/genblk1[1].mult/added[1] ,
         \lamb/scale_ts0/genblk1[1].mult/added[2] ,
         \lamb/scale_ts0/genblk1[1].mult/added[3] ,
         \lamb/scale_ts0/genblk1[1].mult/added[4] ,
         \lamb/scale_ts0/genblk1[1].mult/logA[0] ,
         \lamb/scale_ts0/genblk1[1].mult/logA[1] ,
         \lamb/scale_ts0/genblk1[1].mult/logA[2] ,
         \lamb/scale_ts0/genblk1[1].mult/logA[3] ,
         \lamb/scale_ts0/genblk1[0].mult/added[1] ,
         \lamb/scale_ts0/genblk1[0].mult/added[2] ,
         \lamb/scale_ts0/genblk1[0].mult/added[3] ,
         \lamb/scale_ts0/genblk1[0].mult/added[4] ,
         \lamb/scale_ts0/genblk1[0].mult/logA[0] ,
         \lamb/scale_ts0/genblk1[0].mult/logA[1] ,
         \lamb/scale_ts0/genblk1[0].mult/logA[2] ,
         \lamb/scale_ts0/genblk1[0].mult/logA[3] , \add_x_79/n4 ,
         \add_x_79/n3 , \add_x_79/n2 , \add_x_79/n1 , \add_x_78/n4 ,
         \add_x_78/n3 , \add_x_78/n2 , \add_x_78/n1 , \add_x_77/n4 ,
         \add_x_77/n3 , \add_x_77/n2 , \add_x_77/n1 , \add_x_73/n4 ,
         \add_x_73/n3 , \add_x_73/n2 , \add_x_73/n1 , \add_x_72/n4 ,
         \add_x_72/n3 , \add_x_72/n2 , \add_x_72/n1 , \add_x_71/n4 ,
         \add_x_71/n3 , \add_x_71/n2 , \add_x_71/n1 , \add_x_70/n4 ,
         \add_x_70/n3 , \add_x_70/n2 , \add_x_70/n1 , \add_x_69/n4 ,
         \add_x_69/n3 , \add_x_69/n2 , \add_x_69/n1 , \add_x_68/n4 ,
         \add_x_68/n3 , \add_x_68/n2 , \add_x_68/n1 , \add_x_67/n4 ,
         \add_x_67/n3 , \add_x_67/n2 , \add_x_67/n1 , \add_x_66/n4 ,
         \add_x_66/n3 , \add_x_66/n2 , \add_x_66/n1 , \add_x_65/n4 ,
         \add_x_65/n3 , \add_x_65/n2 , \add_x_65/n1 , \add_x_64/n4 ,
         \add_x_64/n3 , \add_x_64/n2 , \add_x_64/n1 , \add_x_63/n4 ,
         \add_x_63/n3 , \add_x_63/n2 , \add_x_63/n1 , \add_x_60/n4 ,
         \add_x_60/n3 , \add_x_60/n2 , \add_x_60/n1 , \add_x_59/n4 ,
         \add_x_59/n3 , \add_x_59/n2 , \add_x_59/n1 , \add_x_58/n4 ,
         \add_x_58/n3 , \add_x_58/n2 , \add_x_58/n1 , \add_x_56/n4 ,
         \add_x_56/n3 , \add_x_56/n2 , \add_x_56/n1 , \add_x_55/n4 ,
         \add_x_55/n3 , \add_x_55/n2 , \add_x_55/n1 , \add_x_54/n4 ,
         \add_x_54/n3 , \add_x_54/n2 , \add_x_54/n1 , \add_x_53/n4 ,
         \add_x_53/n3 , \add_x_53/n2 , \add_x_53/n1 , \add_x_52/n4 ,
         \add_x_52/n3 , \add_x_52/n2 , \add_x_52/n1 , \add_x_51/n4 ,
         \add_x_51/n3 , \add_x_51/n2 , \add_x_51/n1 , \add_x_50/n4 ,
         \add_x_50/n3 , \add_x_50/n2 , \add_x_50/n1 , \add_x_49/n4 ,
         \add_x_49/n3 , \add_x_49/n2 , \add_x_49/n1 , \add_x_46/n4 ,
         \add_x_46/n3 , \add_x_46/n2 , \add_x_46/n1 , \add_x_45/n4 ,
         \add_x_45/n3 , \add_x_45/n2 , \add_x_45/n1 , \add_x_42/n4 ,
         \add_x_42/n3 , \add_x_42/n2 , \add_x_42/n1 , \add_x_41/n4 ,
         \add_x_41/n3 , \add_x_41/n2 , \add_x_41/n1 , n9905, n9906, n9907,
         n9909, n9911, n9912, n9913, n9917, n16299, n16300, n16301, n16302,
         n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310,
         n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318,
         n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326,
         n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334,
         n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342,
         n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350,
         n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358,
         n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366,
         n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374,
         n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382,
         n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390,
         n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398,
         n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406,
         n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414,
         n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422,
         n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430,
         n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438,
         n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446,
         n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454,
         n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462,
         n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470,
         n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478,
         n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486,
         n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494,
         n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502,
         n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510,
         n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518,
         n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526,
         n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534,
         n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542,
         n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550,
         n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558,
         n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566,
         n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574,
         n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582,
         n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590,
         n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598,
         n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606,
         n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614,
         n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622,
         n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630,
         n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638,
         n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646,
         n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654,
         n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662,
         n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670,
         n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678,
         n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686,
         n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694,
         n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702,
         n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710,
         n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718,
         n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726,
         n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734,
         n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742,
         n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750,
         n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758,
         n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766,
         n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774,
         n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782,
         n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790,
         n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798,
         n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806,
         n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814,
         n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822,
         n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830,
         n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838,
         n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846,
         n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854,
         n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862,
         n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870,
         n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878,
         n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886,
         n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894,
         n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902,
         n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910,
         n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918,
         n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926,
         n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934,
         n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942,
         n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950,
         n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958,
         n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966,
         n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974,
         n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982,
         n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990,
         n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998,
         n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006,
         n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014,
         n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022,
         n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030,
         n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038,
         n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046,
         n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054,
         n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062,
         n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070,
         n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078,
         n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086,
         n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094,
         n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102,
         n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110,
         n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118,
         n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126,
         n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134,
         n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142,
         n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150,
         n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158,
         n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166,
         n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174,
         n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182,
         n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190,
         n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198,
         n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206,
         n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214,
         n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222,
         n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230,
         n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238,
         n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246,
         n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254,
         n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262,
         n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270,
         n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278,
         n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286,
         n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294,
         n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302,
         n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310,
         n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318,
         n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326,
         n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334,
         n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342,
         n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350,
         n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358,
         n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366,
         n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374,
         n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382,
         n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390,
         n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398,
         n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406,
         n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414,
         n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422,
         n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430,
         n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438,
         n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446,
         n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454,
         n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462,
         n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470,
         n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478,
         n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486,
         n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494,
         n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502,
         n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510,
         n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518,
         n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526,
         n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534,
         n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542,
         n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550,
         n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558,
         n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566,
         n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574,
         n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582,
         n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590,
         n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598,
         n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606,
         n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614,
         n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622,
         n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630,
         n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638,
         n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646,
         n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654,
         n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662,
         n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670,
         n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678,
         n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686,
         n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694,
         n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702,
         n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710,
         n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718,
         n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726,
         n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734,
         n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742,
         n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750,
         n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758,
         n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766,
         n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774,
         n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782,
         n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790,
         n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798,
         n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806,
         n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814,
         n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822,
         n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830,
         n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838,
         n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846,
         n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854,
         n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862,
         n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870,
         n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878,
         n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886,
         n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894,
         n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902,
         n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910,
         n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
         n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926,
         n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934,
         n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942,
         n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950,
         n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958,
         n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966,
         n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974,
         n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982,
         n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990,
         n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998,
         n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006,
         n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014,
         n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022,
         n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030,
         n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038,
         n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046,
         n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054,
         n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062,
         n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070,
         n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078,
         n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086,
         n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094,
         n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102,
         n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110,
         n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118,
         n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126,
         n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134,
         n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142,
         n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150,
         n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158,
         n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166,
         n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174,
         n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182,
         n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190,
         n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198,
         n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206,
         n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214,
         n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222,
         n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230,
         n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238,
         n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246,
         n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254,
         n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262,
         n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270,
         n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278,
         n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286,
         n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294,
         n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302,
         n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310,
         n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318,
         n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326,
         n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334,
         n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342,
         n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350,
         n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358,
         n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366,
         n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374,
         n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382,
         n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390,
         n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398,
         n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406,
         n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414,
         n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422,
         n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430,
         n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438,
         n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446,
         n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454,
         n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462,
         n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470,
         n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478,
         n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486,
         n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494,
         n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502,
         n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510,
         n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518,
         n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526,
         n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534,
         n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542,
         n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550,
         n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558,
         n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566,
         n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574,
         n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582,
         n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590,
         n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598,
         n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606,
         n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614,
         n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622,
         n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630,
         n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638,
         n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646,
         n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654,
         n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662,
         n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670,
         n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678,
         n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686,
         n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694,
         n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702,
         n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710,
         n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718,
         n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726,
         n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734,
         n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742,
         n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750,
         n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758,
         n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766,
         n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774,
         n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782,
         n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790,
         n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798,
         n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806,
         n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814,
         n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822,
         n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830,
         n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838,
         n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846,
         n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854,
         n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862,
         n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870,
         n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878,
         n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886,
         n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894,
         n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902,
         n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910,
         n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918,
         n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926,
         n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934,
         n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942,
         n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950,
         n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958,
         n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966,
         n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974,
         n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982,
         n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990,
         n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998,
         n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006,
         n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014,
         n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022,
         n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030,
         n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038,
         n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046,
         n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054,
         n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062,
         n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070,
         n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078,
         n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086,
         n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094,
         n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102,
         n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110,
         n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118,
         n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126,
         n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134,
         n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142,
         n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150,
         n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158,
         n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166,
         n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174,
         n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182,
         n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190,
         n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198,
         n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206,
         n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214,
         n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222,
         n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230,
         n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238,
         n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246,
         n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254,
         n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262,
         n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270,
         n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278,
         n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286,
         n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294,
         n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302,
         n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310,
         n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318,
         n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326,
         n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334,
         n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342,
         n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350,
         n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358,
         n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366,
         n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374,
         n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382,
         n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390,
         n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398,
         n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406,
         n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414,
         n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422,
         n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430,
         n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438,
         n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446,
         n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454,
         n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462,
         n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470,
         n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478,
         n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486,
         n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494,
         n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502,
         n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510,
         n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518,
         n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526,
         n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534,
         n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542,
         n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550,
         n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558,
         n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566,
         n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574,
         n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582,
         n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590,
         n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598,
         n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606,
         n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614,
         n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622,
         n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630,
         n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638,
         n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646,
         n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654,
         n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662,
         n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670,
         n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678,
         n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686,
         n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694,
         n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702,
         n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710,
         n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718,
         n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726,
         n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734,
         n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742,
         n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750,
         n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758,
         n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766,
         n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774,
         n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782;

  HAX1 \add_x_79/U5  ( .A(n16781), .B(\lamb/scale_ts0/genblk1[0].mult/logA[3] ), .YC(\add_x_79/n4 ), .YS(\lamb/scale_ts0/genblk1[0].mult/added[4] ) );
  FAX1 \add_x_79/U4  ( .A(n17124), .B(n16710), .C(\add_x_79/n4 ), .YC(
        \add_x_79/n3 ), .YS(\lamb/scale_ts0/genblk1[0].mult/added[3] ) );
  FAX1 \add_x_79/U3  ( .A(n16314), .B(n17028), .C(\add_x_79/n3 ), .YC(
        \add_x_79/n2 ), .YS(\lamb/scale_ts0/genblk1[0].mult/added[2] ) );
  FAX1 \add_x_79/U2  ( .A(n16316), .B(\lamb/scale_ts0/genblk1[0].mult/logA[0] ), .C(\add_x_79/n2 ), .YC(\add_x_79/n1 ), .YS(
        \lamb/scale_ts0/genblk1[0].mult/added[1] ) );
  HAX1 \add_x_78/U5  ( .A(n16781), .B(\lamb/scale_ts0/genblk1[1].mult/logA[3] ), .YC(\add_x_78/n4 ), .YS(\lamb/scale_ts0/genblk1[1].mult/added[4] ) );
  FAX1 \add_x_78/U4  ( .A(n17124), .B(n16673), .C(\add_x_78/n4 ), .YC(
        \add_x_78/n3 ), .YS(\lamb/scale_ts0/genblk1[1].mult/added[3] ) );
  FAX1 \add_x_78/U3  ( .A(n16314), .B(n16695), .C(\add_x_78/n3 ), .YC(
        \add_x_78/n2 ), .YS(\lamb/scale_ts0/genblk1[1].mult/added[2] ) );
  FAX1 \add_x_78/U2  ( .A(n16316), .B(\lamb/scale_ts0/genblk1[1].mult/logA[0] ), .C(\add_x_78/n2 ), .YC(\add_x_78/n1 ), .YS(
        \lamb/scale_ts0/genblk1[1].mult/added[1] ) );
  HAX1 \add_x_77/U5  ( .A(n16781), .B(\lamb/scale_ts0/genblk1[2].mult/logA[3] ), .YC(\add_x_77/n4 ), .YS(\lamb/scale_ts0/genblk1[2].mult/added[4] ) );
  FAX1 \add_x_77/U4  ( .A(n17124), .B(n16709), .C(\add_x_77/n4 ), .YC(
        \add_x_77/n3 ), .YS(\lamb/scale_ts0/genblk1[2].mult/added[3] ) );
  FAX1 \add_x_77/U3  ( .A(n16314), .B(n17068), .C(\add_x_77/n3 ), .YC(
        \add_x_77/n2 ), .YS(\lamb/scale_ts0/genblk1[2].mult/added[2] ) );
  FAX1 \add_x_77/U2  ( .A(n16316), .B(\lamb/scale_ts0/genblk1[2].mult/logA[0] ), .C(\add_x_77/n2 ), .YC(\add_x_77/n1 ), .YS(
        \lamb/scale_ts0/genblk1[2].mult/added[1] ) );
  HAX1 \add_x_73/U5  ( .A(n16781), .B(\lamb/scale_ds1/genblk1[1].mult/logA[3] ), .YC(\add_x_73/n4 ), .YS(\lamb/scale_ds1/genblk1[1].mult/added[4] ) );
  FAX1 \add_x_73/U4  ( .A(n17124), .B(\lamb/scale_ds1/genblk1[1].mult/logA[2] ), .C(\add_x_73/n4 ), .YC(\add_x_73/n3 ), .YS(
        \lamb/scale_ds1/genblk1[1].mult/added[3] ) );
  FAX1 \add_x_73/U3  ( .A(n16314), .B(n16672), .C(\add_x_73/n3 ), .YC(
        \add_x_73/n2 ), .YS(\lamb/scale_ds1/genblk1[1].mult/added[2] ) );
  FAX1 \add_x_73/U2  ( .A(n16316), .B(n16699), .C(\add_x_73/n2 ), .YC(
        \add_x_73/n1 ), .YS(\lamb/scale_ds1/genblk1[1].mult/added[1] ) );
  HAX1 \add_x_72/U5  ( .A(n16781), .B(\lamb/scale_ds1/genblk1[2].mult/logA[3] ), .YC(\add_x_72/n4 ), .YS(\lamb/scale_ds1/genblk1[2].mult/added[4] ) );
  FAX1 \add_x_72/U4  ( .A(n17124), .B(n9905), .C(\add_x_72/n4 ), .YC(
        \add_x_72/n3 ), .YS(\lamb/scale_ds1/genblk1[2].mult/added[3] ) );
  FAX1 \add_x_72/U3  ( .A(n16314), .B(n16701), .C(\add_x_72/n3 ), .YC(
        \add_x_72/n2 ), .YS(\lamb/scale_ds1/genblk1[2].mult/added[2] ) );
  FAX1 \add_x_72/U2  ( .A(n16316), .B(\lamb/scale_ds1/genblk1[2].mult/logA[0] ), .C(\add_x_72/n2 ), .YC(\add_x_72/n1 ), .YS(
        \lamb/scale_ds1/genblk1[2].mult/added[1] ) );
  HAX1 \add_x_71/U5  ( .A(n16781), .B(\lamb/scale_ds1/genblk1[3].mult/logA[3] ), .YC(\add_x_71/n4 ), .YS(\lamb/scale_ds1/genblk1[3].mult/added[4] ) );
  FAX1 \add_x_71/U4  ( .A(n17124), .B(\lamb/scale_ds1/genblk1[3].mult/logA[2] ), .C(\add_x_71/n4 ), .YC(\add_x_71/n3 ), .YS(
        \lamb/scale_ds1/genblk1[3].mult/added[3] ) );
  FAX1 \add_x_71/U3  ( .A(n16314), .B(n9912), .C(\add_x_71/n3 ), .YC(
        \add_x_71/n2 ), .YS(\lamb/scale_ds1/genblk1[3].mult/added[2] ) );
  FAX1 \add_x_71/U2  ( .A(n16316), .B(n9911), .C(\add_x_71/n2 ), .YC(
        \add_x_71/n1 ), .YS(\lamb/scale_ds1/genblk1[3].mult/added[1] ) );
  HAX1 \add_x_70/U5  ( .A(\lamb/scale_ts1/genblk1[0].mult/logB[3] ), .B(
        \lamb/scale_ts1/genblk1[0].mult/logA[3] ), .YC(\add_x_70/n4 ), .YS(
        \lamb/scale_ts1/genblk1[0].mult/added[4] ) );
  FAX1 \add_x_70/U4  ( .A(n17106), .B(\lamb/scale_ts1/genblk1[0].mult/logA[2] ), .C(\add_x_70/n4 ), .YC(\add_x_70/n3 ), .YS(
        \lamb/scale_ts1/genblk1[0].mult/added[3] ) );
  FAX1 \add_x_70/U3  ( .A(n16776), .B(\lamb/scale_ts1/genblk1[0].mult/logA[1] ), .C(\add_x_70/n3 ), .YC(\add_x_70/n2 ), .YS(
        \lamb/scale_ts1/genblk1[0].mult/added[2] ) );
  FAX1 \add_x_70/U2  ( .A(\lamb/scale_ts1/genblk1[0].mult/logB[0] ), .B(
        \lamb/scale_ts1/genblk1[0].mult/logA[0] ), .C(\add_x_70/n2 ), .YC(
        \add_x_70/n1 ), .YS(\lamb/scale_ts1/genblk1[0].mult/added[1] ) );
  HAX1 \add_x_69/U5  ( .A(\lamb/scale_ts1/genblk1[0].mult/logB[3] ), .B(
        \lamb/scale_ts1/genblk1[1].mult/logA[3] ), .YC(\add_x_69/n4 ), .YS(
        \lamb/scale_ts1/genblk1[1].mult/added[4] ) );
  FAX1 \add_x_69/U4  ( .A(n17106), .B(n16700), .C(\add_x_69/n4 ), .YC(
        \add_x_69/n3 ), .YS(\lamb/scale_ts1/genblk1[1].mult/added[3] ) );
  FAX1 \add_x_69/U3  ( .A(n16776), .B(n16671), .C(\add_x_69/n3 ), .YC(
        \add_x_69/n2 ), .YS(\lamb/scale_ts1/genblk1[1].mult/added[2] ) );
  FAX1 \add_x_69/U2  ( .A(\lamb/scale_ts1/genblk1[0].mult/logB[0] ), .B(n16310), .C(\add_x_69/n2 ), .YC(\add_x_69/n1 ), .YS(
        \lamb/scale_ts1/genblk1[1].mult/added[1] ) );
  HAX1 \add_x_68/U5  ( .A(\lamb/scale_ts1/genblk1[0].mult/logB[3] ), .B(n16305), .YC(\add_x_68/n4 ), .YS(\lamb/scale_ts1/genblk1[2].mult/added[4] ) );
  FAX1 \add_x_68/U4  ( .A(n17106), .B(n16694), .C(\add_x_68/n4 ), .YC(
        \add_x_68/n3 ), .YS(\lamb/scale_ts1/genblk1[2].mult/added[3] ) );
  FAX1 \add_x_68/U3  ( .A(n16776), .B(\lamb/scale_ts1/genblk1[2].mult/logA[1] ), .C(\add_x_68/n3 ), .YC(\add_x_68/n2 ), .YS(
        \lamb/scale_ts1/genblk1[2].mult/added[2] ) );
  FAX1 \add_x_68/U2  ( .A(\lamb/scale_ts1/genblk1[0].mult/logB[0] ), .B(
        \lamb/scale_ts1/genblk1[2].mult/logA[0] ), .C(\add_x_68/n2 ), .YC(
        \add_x_68/n1 ), .YS(\lamb/scale_ts1/genblk1[2].mult/added[1] ) );
  HAX1 \add_x_67/U5  ( .A(\lamb/scale_ts1/genblk1[0].mult/logB[3] ), .B(n17031), .YC(\add_x_67/n4 ), .YS(\lamb/scale_ts1/genblk1[3].mult/added[4] ) );
  FAX1 \add_x_67/U4  ( .A(n17106), .B(\lamb/scale_ls2/genblk1[1].mult/logA[2] ), .C(\add_x_67/n4 ), .YC(\add_x_67/n3 ), .YS(
        \lamb/scale_ts1/genblk1[3].mult/added[3] ) );
  FAX1 \add_x_67/U3  ( .A(n16776), .B(\lamb/scale_ts1/genblk1[3].mult/logA[1] ), .C(\add_x_67/n3 ), .YC(\add_x_67/n2 ), .YS(
        \lamb/scale_ts1/genblk1[3].mult/added[2] ) );
  FAX1 \add_x_67/U2  ( .A(\lamb/scale_ts1/genblk1[0].mult/logB[0] ), .B(
        \lamb/scale_ts1/genblk1[3].mult/logA[0] ), .C(\add_x_67/n2 ), .YC(
        \add_x_67/n1 ), .YS(\lamb/scale_ts1/genblk1[3].mult/added[1] ) );
  HAX1 \add_x_66/U5  ( .A(n16770), .B(\lamb/scale_ls2/genblk1[0].mult/logA[3] ), .YC(\add_x_66/n4 ), .YS(\lamb/scale_ls2/genblk1[0].mult/added[4] ) );
  FAX1 \add_x_66/U4  ( .A(n16782), .B(n16693), .C(\add_x_66/n4 ), .YC(
        \add_x_66/n3 ), .YS(\lamb/scale_ls2/genblk1[0].mult/added[3] ) );
  FAX1 \add_x_66/U3  ( .A(n17117), .B(\lamb/scale_ls2/genblk1[0].mult/logA[1] ), .C(\add_x_66/n3 ), .YC(\add_x_66/n2 ), .YS(
        \lamb/scale_ls2/genblk1[0].mult/added[2] ) );
  FAX1 \add_x_66/U2  ( .A(\lamb/scale_ls2/genblk1[0].mult/logB[0] ), .B(
        \lamb/scale_ls2/genblk1[0].mult/logA[0] ), .C(\add_x_66/n2 ), .YC(
        \add_x_66/n1 ), .YS(\lamb/scale_ls2/genblk1[0].mult/added[1] ) );
  HAX1 \add_x_65/U5  ( .A(n16770), .B(n17031), .YC(\add_x_65/n4 ), .YS(
        \lamb/scale_ls2/genblk1[1].mult/added[4] ) );
  FAX1 \add_x_65/U4  ( .A(n16782), .B(\lamb/scale_ls2/genblk1[1].mult/logA[2] ), .C(\add_x_65/n4 ), .YC(\add_x_65/n3 ), .YS(
        \lamb/scale_ls2/genblk1[1].mult/added[3] ) );
  FAX1 \add_x_65/U3  ( .A(n17117), .B(\lamb/scale_ts1/genblk1[3].mult/logA[1] ), .C(\add_x_65/n3 ), .YC(\add_x_65/n2 ), .YS(
        \lamb/scale_ls2/genblk1[1].mult/added[2] ) );
  FAX1 \add_x_65/U2  ( .A(\lamb/scale_ls2/genblk1[0].mult/logB[0] ), .B(
        \lamb/scale_ts1/genblk1[3].mult/logA[0] ), .C(\add_x_65/n2 ), .YC(
        \add_x_65/n1 ), .YS(\lamb/scale_ls2/genblk1[1].mult/added[1] ) );
  HAX1 \add_x_64/U5  ( .A(n16770), .B(n16781), .YC(\add_x_64/n4 ), .YS(
        \lamb/scale_ls2/genblk1[2].mult/added[4] ) );
  FAX1 \add_x_64/U4  ( .A(n16782), .B(n17124), .C(\add_x_64/n4 ), .YC(
        \add_x_64/n3 ), .YS(\lamb/scale_ls2/genblk1[2].mult/added[3] ) );
  FAX1 \add_x_64/U3  ( .A(n17117), .B(n16314), .C(\add_x_64/n3 ), .YC(
        \add_x_64/n2 ), .YS(\lamb/scale_ls2/genblk1[2].mult/added[2] ) );
  FAX1 \add_x_64/U2  ( .A(\lamb/scale_ls2/genblk1[0].mult/logB[0] ), .B(n16316), .C(\add_x_64/n2 ), .YC(\add_x_64/n1 ), .YS(
        \lamb/scale_ls2/genblk1[2].mult/added[1] ) );
  HAX1 \add_x_63/U5  ( .A(n17085), .B(\lamb/scale_bs2/genblk1[0].mult/logA[3] ), .YC(\add_x_63/n4 ), .YS(\lamb/scale_bs2/genblk1[0].mult/added[4] ) );
  FAX1 \add_x_63/U4  ( .A(\lamb/scale_bs2/genblk1[1].mult/added[3] ), .B(
        \lamb/scale_bs2/genblk1[0].mult/logA[2] ), .C(\add_x_63/n4 ), .YC(
        \add_x_63/n3 ), .YS(\lamb/scale_bs2/genblk1[0].mult/added[3] ) );
  FAX1 \add_x_63/U3  ( .A(n17105), .B(n16315), .C(\add_x_63/n3 ), .YC(
        \add_x_63/n2 ), .YS(\lamb/scale_bs2/genblk1[0].mult/added[2] ) );
  FAX1 \add_x_63/U2  ( .A(n16301), .B(\lamb/scale_bs2/genblk1[0].mult/logA[0] ), .C(\add_x_63/n2 ), .YC(\add_x_63/n1 ), .YS(
        \lamb/scale_bs2/genblk1[0].mult/added[1] ) );
  HAX1 \add_x_60/U5  ( .A(n16770), .B(\lamb/scale_ds2/genblk1[1].mult/logA[3] ), .YC(\add_x_60/n4 ), .YS(\lamb/scale_ds2/genblk1[1].mult/added[4] ) );
  FAX1 \add_x_60/U4  ( .A(n16782), .B(n16925), .C(\add_x_60/n4 ), .YC(
        \add_x_60/n3 ), .YS(\lamb/scale_ds2/genblk1[1].mult/added[3] ) );
  FAX1 \add_x_60/U3  ( .A(n17117), .B(n16692), .C(\add_x_60/n3 ), .YC(
        \add_x_60/n2 ), .YS(\lamb/scale_ds2/genblk1[1].mult/added[2] ) );
  FAX1 \add_x_60/U2  ( .A(\lamb/scale_ls2/genblk1[0].mult/logB[0] ), .B(
        \lamb/scale_ds2/genblk1[1].mult/logA[0] ), .C(\add_x_60/n2 ), .YC(
        \add_x_60/n1 ), .YS(\lamb/scale_ds2/genblk1[1].mult/added[1] ) );
  HAX1 \add_x_59/U5  ( .A(n16770), .B(n16860), .YC(\add_x_59/n4 ), .YS(
        \lamb/scale_ds2/genblk1[2].mult/added[4] ) );
  FAX1 \add_x_59/U4  ( .A(n16782), .B(n16691), .C(\add_x_59/n4 ), .YC(
        \add_x_59/n3 ), .YS(\lamb/scale_ds2/genblk1[2].mult/added[3] ) );
  FAX1 \add_x_59/U3  ( .A(n17117), .B(n16690), .C(\add_x_59/n3 ), .YC(
        \add_x_59/n2 ), .YS(\lamb/scale_ds2/genblk1[2].mult/added[2] ) );
  FAX1 \add_x_59/U2  ( .A(\lamb/scale_ls2/genblk1[0].mult/logB[0] ), .B(
        \lamb/scale_ds2/genblk1[2].mult/logA[0] ), .C(\add_x_59/n2 ), .YC(
        \add_x_59/n1 ), .YS(\lamb/scale_ds2/genblk1[2].mult/added[1] ) );
  HAX1 \add_x_58/U5  ( .A(n16770), .B(\lamb/scale_ds2/genblk1[3].mult/logA[3] ), .YC(\add_x_58/n4 ), .YS(\lamb/scale_ds2/genblk1[3].mult/added[4] ) );
  FAX1 \add_x_58/U4  ( .A(n16782), .B(n16698), .C(\add_x_58/n4 ), .YC(
        \add_x_58/n3 ), .YS(\lamb/scale_ds2/genblk1[3].mult/added[3] ) );
  FAX1 \add_x_58/U3  ( .A(n17117), .B(n16689), .C(\add_x_58/n3 ), .YC(
        \add_x_58/n2 ), .YS(\lamb/scale_ds2/genblk1[3].mult/added[2] ) );
  FAX1 \add_x_58/U2  ( .A(\lamb/scale_ls2/genblk1[0].mult/logB[0] ), .B(
        \lamb/scale_ds2/genblk1[3].mult/logA[0] ), .C(\add_x_58/n2 ), .YC(
        \add_x_58/n1 ), .YS(\lamb/scale_ds2/genblk1[3].mult/added[1] ) );
  HAX1 \add_x_56/U5  ( .A(n17085), .B(\lamb/scale_ts2/genblk1[1].mult/logA[3] ), .YC(\add_x_56/n4 ), .YS(\lamb/scale_ts2/genblk1[1].mult/added[4] ) );
  FAX1 \add_x_56/U4  ( .A(\lamb/scale_bs2/genblk1[1].mult/added[3] ), .B(
        n16688), .C(\add_x_56/n4 ), .YC(\add_x_56/n3 ), .YS(
        \lamb/scale_ts2/genblk1[1].mult/added[3] ) );
  FAX1 \add_x_56/U3  ( .A(n17105), .B(n16677), .C(\add_x_56/n3 ), .YC(
        \add_x_56/n2 ), .YS(\lamb/scale_ts2/genblk1[1].mult/added[2] ) );
  FAX1 \add_x_56/U2  ( .A(n16301), .B(\lamb/scale_ts2/genblk1[1].mult/logA[0] ), .C(\add_x_56/n2 ), .YC(\add_x_56/n1 ), .YS(
        \lamb/scale_ts2/genblk1[1].mult/added[1] ) );
  HAX1 \add_x_55/U5  ( .A(n17085), .B(\lamb/scale_ts2/genblk1[2].mult/logA[3] ), .YC(\add_x_55/n4 ), .YS(\lamb/scale_ts2/genblk1[2].mult/added[4] ) );
  FAX1 \add_x_55/U4  ( .A(\lamb/scale_bs2/genblk1[1].mult/added[3] ), .B(
        \lamb/scale_ts2/genblk1[2].mult/logA[2] ), .C(\add_x_55/n4 ), .YC(
        \add_x_55/n3 ), .YS(\lamb/scale_ts2/genblk1[2].mult/added[3] ) );
  FAX1 \add_x_55/U3  ( .A(n17105), .B(n16687), .C(\add_x_55/n3 ), .YC(
        \add_x_55/n2 ), .YS(\lamb/scale_ts2/genblk1[2].mult/added[2] ) );
  FAX1 \add_x_55/U2  ( .A(n16301), .B(n9906), .C(\add_x_55/n2 ), .YC(
        \add_x_55/n1 ), .YS(\lamb/scale_ts2/genblk1[2].mult/added[1] ) );
  HAX1 \add_x_54/U5  ( .A(n17085), .B(\lamb/scale_ts2/genblk1[3].mult/logA[3] ), .YC(\add_x_54/n4 ), .YS(\lamb/scale_ts2/genblk1[3].mult/added[4] ) );
  FAX1 \add_x_54/U4  ( .A(\lamb/scale_bs2/genblk1[1].mult/added[3] ), .B(
        \lamb/scale_ts2/genblk1[3].mult/logA[2] ), .C(\add_x_54/n4 ), .YC(
        \add_x_54/n3 ), .YS(\lamb/scale_ts2/genblk1[3].mult/added[3] ) );
  FAX1 \add_x_54/U3  ( .A(n17105), .B(n16686), .C(\add_x_54/n3 ), .YC(
        \add_x_54/n2 ), .YS(\lamb/scale_ts2/genblk1[3].mult/added[2] ) );
  FAX1 \add_x_54/U2  ( .A(n16301), .B(n9913), .C(\add_x_54/n2 ), .YC(
        \add_x_54/n1 ), .YS(\lamb/scale_ts2/genblk1[3].mult/added[1] ) );
  HAX1 \add_x_53/U5  ( .A(\lamb/scale_ls3/genblk1[0].mult/logB[3] ), .B(
        \lamb/scale_ls3/genblk1[0].mult/logA[3] ), .YC(\add_x_53/n4 ), .YS(
        \lamb/scale_ls3/genblk1[0].mult/added[4] ) );
  FAX1 \add_x_53/U4  ( .A(n17109), .B(n16685), .C(\add_x_53/n4 ), .YC(
        \add_x_53/n3 ), .YS(\lamb/scale_ls3/genblk1[0].mult/added[3] ) );
  FAX1 \add_x_53/U3  ( .A(n16777), .B(n16684), .C(\add_x_53/n3 ), .YC(
        \add_x_53/n2 ), .YS(\lamb/scale_ls3/genblk1[0].mult/added[2] ) );
  FAX1 \add_x_53/U2  ( .A(n16302), .B(n16300), .C(\add_x_53/n2 ), .YC(
        \add_x_53/n1 ), .YS(\lamb/scale_ls3/genblk1[0].mult/added[1] ) );
  HAX1 \add_x_52/U5  ( .A(\lamb/scale_ls3/genblk1[0].mult/logB[3] ), .B(
        \lamb/scale_ls3/genblk1[1].mult/logA[3] ), .YC(\add_x_52/n4 ), .YS(
        \lamb/scale_ls3/genblk1[1].mult/added[4] ) );
  FAX1 \add_x_52/U4  ( .A(n17109), .B(n16670), .C(\add_x_52/n4 ), .YC(
        \add_x_52/n3 ), .YS(\lamb/scale_ls3/genblk1[1].mult/added[3] ) );
  FAX1 \add_x_52/U3  ( .A(n16777), .B(n16683), .C(\add_x_52/n3 ), .YC(
        \add_x_52/n2 ), .YS(\lamb/scale_ls3/genblk1[1].mult/added[2] ) );
  FAX1 \add_x_52/U2  ( .A(n16302), .B(\lamb/scale_ls3/genblk1[1].mult/logA[0] ), .C(\add_x_52/n2 ), .YC(\add_x_52/n1 ), .YS(
        \lamb/scale_ls3/genblk1[1].mult/added[1] ) );
  HAX1 \add_x_51/U5  ( .A(\lamb/scale_ls3/genblk1[0].mult/logB[3] ), .B(
        \lamb/scale_ls3/genblk1[2].mult/logA[3] ), .YC(\add_x_51/n4 ), .YS(
        \lamb/scale_ls3/genblk1[2].mult/added[4] ) );
  FAX1 \add_x_51/U4  ( .A(n17109), .B(\lamb/scale_ls3/genblk1[2].mult/logA[2] ), .C(\add_x_51/n4 ), .YC(\add_x_51/n3 ), .YS(
        \lamb/scale_ls3/genblk1[2].mult/added[3] ) );
  FAX1 \add_x_51/U3  ( .A(n16777), .B(n16923), .C(\add_x_51/n3 ), .YC(
        \add_x_51/n2 ), .YS(\lamb/scale_ls3/genblk1[2].mult/added[2] ) );
  FAX1 \add_x_51/U2  ( .A(n16302), .B(n16682), .C(\add_x_51/n2 ), .YC(
        \add_x_51/n1 ), .YS(\lamb/scale_ls3/genblk1[2].mult/added[1] ) );
  HAX1 \add_x_50/U5  ( .A(n17084), .B(\lamb/scale_bs3/genblk1[0].mult/logA[3] ), .YC(\add_x_50/n4 ), .YS(\lamb/scale_bs3/genblk1[0].mult/added[4] ) );
  FAX1 \add_x_50/U4  ( .A(n16299), .B(\lamb/scale_bs3/genblk1[0].mult/logA[2] ), .C(\add_x_50/n4 ), .YC(\add_x_50/n3 ), .YS(
        \lamb/scale_bs3/genblk1[0].mult/added[3] ) );
  FAX1 \add_x_50/U3  ( .A(n17104), .B(\lamb/scale_bs3/genblk1[0].mult/logA[1] ), .C(\add_x_50/n3 ), .YC(\add_x_50/n2 ), .YS(
        \lamb/scale_bs3/genblk1[0].mult/added[2] ) );
  FAX1 \add_x_50/U2  ( .A(\lamb/scale_bs3/genblk1[0].mult/logB[0] ), .B(
        \lamb/scale_bs3/genblk1[0].mult/logA[0] ), .C(\add_x_50/n2 ), .YC(
        \add_x_50/n1 ), .YS(\lamb/scale_bs3/genblk1[0].mult/added[1] ) );
  HAX1 \add_x_49/U5  ( .A(n17084), .B(\lamb/scale_bs3/genblk1[1].mult/logA[3] ), .YC(\add_x_49/n4 ), .YS(\lamb/scale_bs3/genblk1[1].mult/added[4] ) );
  FAX1 \add_x_49/U4  ( .A(n16299), .B(n9909), .C(\add_x_49/n4 ), .YC(
        \add_x_49/n3 ), .YS(\lamb/scale_bs3/genblk1[1].mult/added[3] ) );
  FAX1 \add_x_49/U3  ( .A(n17104), .B(n16303), .C(\add_x_49/n3 ), .YC(
        \add_x_49/n2 ), .YS(\lamb/scale_bs3/genblk1[1].mult/added[2] ) );
  FAX1 \add_x_49/U2  ( .A(\lamb/scale_bs3/genblk1[0].mult/logB[0] ), .B(
        \lamb/scale_bs3/genblk1[1].mult/logA[0] ), .C(\add_x_49/n2 ), .YC(
        \add_x_49/n1 ), .YS(\lamb/scale_bs3/genblk1[1].mult/added[1] ) );
  HAX1 \add_x_46/U5  ( .A(\lamb/scale_ls3/genblk1[0].mult/logB[3] ), .B(
        \lamb/scale_ds3/genblk1[2].mult/logA[3] ), .YC(\add_x_46/n4 ), .YS(
        \lamb/scale_ds3/genblk1[2].mult/added[4] ) );
  FAX1 \add_x_46/U4  ( .A(n17109), .B(n16681), .C(\add_x_46/n4 ), .YC(
        \add_x_46/n3 ), .YS(\lamb/scale_ds3/genblk1[2].mult/added[3] ) );
  FAX1 \add_x_46/U3  ( .A(n16777), .B(n16680), .C(\add_x_46/n3 ), .YC(
        \add_x_46/n2 ), .YS(\lamb/scale_ds3/genblk1[2].mult/added[2] ) );
  FAX1 \add_x_46/U2  ( .A(n16302), .B(n9907), .C(\add_x_46/n2 ), .YC(
        \add_x_46/n1 ), .YS(\lamb/scale_ds3/genblk1[2].mult/added[1] ) );
  HAX1 \add_x_45/U5  ( .A(\lamb/scale_ls3/genblk1[0].mult/logB[3] ), .B(n16852), .YC(\add_x_45/n4 ), .YS(\lamb/scale_ds3/genblk1[3].mult/added[4] ) );
  FAX1 \add_x_45/U4  ( .A(n17109), .B(n16679), .C(\add_x_45/n4 ), .YC(
        \add_x_45/n3 ), .YS(\lamb/scale_ds3/genblk1[3].mult/added[3] ) );
  FAX1 \add_x_45/U3  ( .A(n16777), .B(\lamb/scale_ds3/genblk1[3].mult/logA[1] ), .C(\add_x_45/n3 ), .YC(\add_x_45/n2 ), .YS(
        \lamb/scale_ds3/genblk1[3].mult/added[2] ) );
  FAX1 \add_x_45/U2  ( .A(n16302), .B(\lamb/scale_ds3/genblk1[3].mult/logA[0] ), .C(\add_x_45/n2 ), .YC(\add_x_45/n1 ), .YS(
        \lamb/scale_ds3/genblk1[3].mult/added[1] ) );
  HAX1 \add_x_42/U5  ( .A(n17084), .B(\lamb/scale_ts3/genblk1[2].mult/logA[3] ), .YC(\add_x_42/n4 ), .YS(\lamb/scale_ts3/genblk1[2].mult/added[4] ) );
  FAX1 \add_x_42/U4  ( .A(n16299), .B(n16924), .C(\add_x_42/n4 ), .YC(
        \add_x_42/n3 ), .YS(\lamb/scale_ts3/genblk1[2].mult/added[3] ) );
  FAX1 \add_x_42/U3  ( .A(n17104), .B(\lamb/scale_ts3/genblk1[2].mult/logA[1] ), .C(\add_x_42/n3 ), .YC(\add_x_42/n2 ), .YS(
        \lamb/scale_ts3/genblk1[2].mult/added[2] ) );
  FAX1 \add_x_42/U2  ( .A(\lamb/scale_bs3/genblk1[0].mult/logB[0] ), .B(
        \lamb/scale_ts3/genblk1[2].mult/logA[0] ), .C(\add_x_42/n2 ), .YC(
        \add_x_42/n1 ), .YS(\lamb/scale_ts3/genblk1[2].mult/added[1] ) );
  HAX1 \add_x_41/U5  ( .A(n17084), .B(\lamb/scale_ts3/genblk1[3].mult/logA[3] ), .YC(\add_x_41/n4 ), .YS(\lamb/scale_ts3/genblk1[3].mult/added[4] ) );
  FAX1 \add_x_41/U4  ( .A(n16299), .B(n16678), .C(\add_x_41/n4 ), .YC(
        \add_x_41/n3 ), .YS(\lamb/scale_ts3/genblk1[3].mult/added[3] ) );
  FAX1 \add_x_41/U3  ( .A(n17104), .B(\lamb/scale_ts3/genblk1[3].mult/logA[1] ), .C(\add_x_41/n3 ), .YC(\add_x_41/n2 ), .YS(
        \lamb/scale_ts3/genblk1[3].mult/added[2] ) );
  FAX1 \add_x_41/U2  ( .A(\lamb/scale_bs3/genblk1[0].mult/logB[0] ), .B(
        \lamb/scale_ts3/genblk1[3].mult/logA[0] ), .C(\add_x_41/n2 ), .YC(
        \add_x_41/n1 ), .YS(\lamb/scale_ts3/genblk1[3].mult/added[1] ) );
  AND2X1 U9524 ( .A(n19081), .B(n16375), .Y(n19146) );
  OR2X1 U9525 ( .A(n18575), .B(n16361), .Y(n18573) );
  AND2X1 U9526 ( .A(n16324), .B(n17966), .Y(n17989) );
  OR2X1 U9527 ( .A(n17654), .B(n16458), .Y(n17700) );
  AND2X1 U9528 ( .A(n19088), .B(n16656), .Y(n19155) );
  INVX1 U9529 ( .A(n19155), .Y(n16317) );
  OR2X1 U9530 ( .A(n17759), .B(n17042), .Y(n17775) );
  INVX1 U9531 ( .A(n17775), .Y(n16318) );
  BUFX2 U9532 ( .A(n17810), .Y(n16319) );
  AND2X1 U9533 ( .A(n16458), .B(n17654), .Y(n17726) );
  INVX1 U9534 ( .A(n17726), .Y(n16320) );
  AND2X1 U9535 ( .A(\lamb/scale_ts2/genblk1[2].mult/added[2] ), .B(n17873), 
        .Y(n17909) );
  INVX1 U9536 ( .A(n17909), .Y(n16321) );
  AND2X1 U9537 ( .A(n17123), .B(n18122), .Y(n18123) );
  INVX1 U9538 ( .A(n18123), .Y(n16322) );
  AND2X1 U9539 ( .A(n19712), .B(n17123), .Y(n18134) );
  INVX1 U9540 ( .A(n18134), .Y(n16323) );
  OR2X1 U9541 ( .A(\lamb/scale_ds2/genblk1[1].mult/added[4] ), .B(
        \add_x_60/n1 ), .Y(n17952) );
  INVX1 U9542 ( .A(n17952), .Y(n16324) );
  AND2X1 U9543 ( .A(n18406), .B(n18405), .Y(n19777) );
  INVX1 U9544 ( .A(n19777), .Y(n16325) );
  AND2X1 U9545 ( .A(n18507), .B(n18390), .Y(n18536) );
  INVX1 U9546 ( .A(n18536), .Y(n16326) );
  OR2X1 U9547 ( .A(n17426), .B(n16524), .Y(n17452) );
  INVX1 U9548 ( .A(n17452), .Y(n16327) );
  AND2X1 U9549 ( .A(n17631), .B(n16386), .Y(n17508) );
  INVX1 U9550 ( .A(n17508), .Y(n16328) );
  AND2X1 U9551 ( .A(\lamb/scale_ts3/genblk1[3].mult/added[4] ), .B(
        \add_x_41/n1 ), .Y(n19125) );
  INVX1 U9552 ( .A(n19125), .Y(n16329) );
  AND2X2 U9553 ( .A(n18979), .B(n18978), .Y(n19019) );
  INVX1 U9554 ( .A(n19019), .Y(n16330) );
  AND2X1 U9555 ( .A(n19055), .B(n16637), .Y(n19060) );
  INVX1 U9556 ( .A(n19060), .Y(n16331) );
  BUFX2 U9557 ( .A(n17845), .Y(n16332) );
  BUFX2 U9558 ( .A(n18106), .Y(n16333) );
  OR2X1 U9559 ( .A(n17018), .B(n17749), .Y(n17753) );
  INVX1 U9560 ( .A(n17753), .Y(n16334) );
  AND2X1 U9561 ( .A(\lamb/scale_bs3/genblk1[0].mult/added[1] ), .B(
        \lamb/scale_bs3/genblk1[0].mult/added[2] ), .Y(n18563) );
  INVX1 U9562 ( .A(n18563), .Y(n16335) );
  AND2X2 U9563 ( .A(n17023), .B(n19330), .Y(n19343) );
  INVX1 U9564 ( .A(n19343), .Y(n16336) );
  AND2X1 U9565 ( .A(\lamb/scale_ts2/genblk1[1].mult/added[3] ), .B(n17977), 
        .Y(n18002) );
  INVX1 U9566 ( .A(n18002), .Y(n16337) );
  BUFX2 U9567 ( .A(n18748), .Y(n16338) );
  BUFX2 U9568 ( .A(n18136), .Y(n16339) );
  AND2X1 U9569 ( .A(n18381), .B(n17642), .Y(n18386) );
  INVX1 U9570 ( .A(n18386), .Y(n16340) );
  AND2X1 U9571 ( .A(n18159), .B(n17004), .Y(n18165) );
  INVX1 U9572 ( .A(n18165), .Y(n16341) );
  OR2X1 U9573 ( .A(n18993), .B(n18996), .Y(n18992) );
  INVX1 U9574 ( .A(n18992), .Y(n16342) );
  AND2X1 U9575 ( .A(\lamb/scale_ls2/genblk1[0].mult/added[2] ), .B(n17052), 
        .Y(n17547) );
  INVX1 U9576 ( .A(n17547), .Y(n16343) );
  AND2X1 U9577 ( .A(n17603), .B(n16485), .Y(n17393) );
  INVX1 U9578 ( .A(n17393), .Y(n16344) );
  AND2X1 U9579 ( .A(n18259), .B(n18260), .Y(n18256) );
  INVX1 U9580 ( .A(n18256), .Y(n16345) );
  INVX1 U9581 ( .A(n16346), .Y(n19177) );
  INVX1 U9582 ( .A(n19149), .Y(n16347) );
  INVX1 U9583 ( .A(n19150), .Y(n16348) );
  INVX1 U9584 ( .A(n19151), .Y(n16349) );
  NOR2X1 U9585 ( .A(n16349), .B(n16350), .Y(n16346) );
  NOR2X1 U9586 ( .A(n16347), .B(n16348), .Y(n16351) );
  INVX1 U9587 ( .A(n16351), .Y(n16350) );
  BUFX2 U9588 ( .A(n19515), .Y(n16352) );
  AND2X1 U9589 ( .A(n18381), .B(n18384), .Y(n18387) );
  INVX1 U9590 ( .A(n18387), .Y(n16353) );
  AND2X1 U9591 ( .A(\lamb/scale_ds1/genblk1[1].mult/added[1] ), .B(
        \lamb/scale_ds1/genblk1[1].mult/added[2] ), .Y(n17774) );
  INVX1 U9592 ( .A(n17774), .Y(n16354) );
  OR2X2 U9593 ( .A(n19114), .B(n19085), .Y(n19152) );
  INVX1 U9594 ( .A(n19152), .Y(n16355) );
  AND2X2 U9595 ( .A(n19121), .B(n19151), .Y(n19179) );
  INVX1 U9596 ( .A(n19179), .Y(n16356) );
  AND2X2 U9597 ( .A(n19386), .B(n19385), .Y(n19391) );
  INVX1 U9598 ( .A(n19391), .Y(n16357) );
  BUFX2 U9599 ( .A(n19186), .Y(n16358) );
  AND2X1 U9600 ( .A(\lamb/scale_bs3/genblk1[0].mult/added[1] ), .B(n18422), 
        .Y(n18566) );
  INVX1 U9601 ( .A(n18566), .Y(n16359) );
  AND2X1 U9602 ( .A(n17043), .B(n19274), .Y(n19279) );
  INVX1 U9603 ( .A(n19279), .Y(n16360) );
  BUFX2 U9604 ( .A(n18589), .Y(n16361) );
  OR2X1 U9605 ( .A(\lamb/scale_ts2/genblk1[2].mult/added[1] ), .B(n17894), .Y(
        n17871) );
  INVX1 U9606 ( .A(n17871), .Y(n16362) );
  BUFX2 U9607 ( .A(n18238), .Y(n16363) );
  BUFX2 U9608 ( .A(n17696), .Y(n16364) );
  AND2X1 U9609 ( .A(\lamb/scale_ls3/genblk1[0].mult/added[2] ), .B(n18491), 
        .Y(n18552) );
  INVX1 U9610 ( .A(n18552), .Y(n16365) );
  BUFX2 U9611 ( .A(n17298), .Y(n16366) );
  BUFX2 U9612 ( .A(n19207), .Y(n16367) );
  OR2X1 U9613 ( .A(n16758), .B(n16747), .Y(n18972) );
  INVX1 U9614 ( .A(n18972), .Y(n16368) );
  AND2X1 U9615 ( .A(\lamb/scale_ts2/genblk1[2].mult/added[2] ), .B(
        \lamb/scale_ts2/genblk1[2].mult/added[1] ), .Y(n17916) );
  INVX1 U9616 ( .A(n17916), .Y(n16369) );
  AND2X1 U9617 ( .A(n18319), .B(n16482), .Y(n18324) );
  INVX1 U9618 ( .A(n18324), .Y(n16370) );
  AND2X1 U9619 ( .A(n19239), .B(n17005), .Y(n19228) );
  INVX1 U9620 ( .A(n19228), .Y(n16371) );
  BUFX2 U9621 ( .A(n19095), .Y(n16372) );
  BUFX2 U9622 ( .A(n18971), .Y(n16373) );
  AND2X1 U9623 ( .A(\lamb/scale_ds2/genblk1[1].mult/added[2] ), .B(n17985), 
        .Y(n17988) );
  INVX1 U9624 ( .A(n17988), .Y(n16374) );
  OR2X1 U9625 ( .A(n19074), .B(n19075), .Y(n19080) );
  INVX1 U9626 ( .A(n19080), .Y(n16375) );
  BUFX2 U9627 ( .A(n18305), .Y(n16376) );
  BUFX2 U9628 ( .A(n19206), .Y(n16377) );
  BUFX2 U9629 ( .A(n19690), .Y(n16378) );
  BUFX2 U9630 ( .A(n18928), .Y(n16379) );
  AND2X1 U9631 ( .A(n18187), .B(n18186), .Y(n18195) );
  INVX1 U9632 ( .A(n18195), .Y(n16380) );
  AND2X2 U9633 ( .A(n18329), .B(n17695), .Y(n18292) );
  INVX1 U9634 ( .A(n18292), .Y(n16381) );
  AND2X2 U9635 ( .A(n18824), .B(n18819), .Y(n18833) );
  AND2X2 U9636 ( .A(n19173), .B(n19196), .Y(n19174) );
  AND2X2 U9637 ( .A(n17744), .B(n17740), .Y(n17747) );
  AND2X2 U9638 ( .A(n18415), .B(n18970), .Y(n18565) );
  AND2X2 U9639 ( .A(n18414), .B(n18970), .Y(n18531) );
  AND2X2 U9640 ( .A(n16361), .B(n18581), .Y(n18720) );
  INVX1 U9641 ( .A(n16384), .Y(n16382) );
  INVX1 U9642 ( .A(n16382), .Y(n16383) );
  AND2X1 U9643 ( .A(n17630), .B(n16576), .Y(n17780) );
  INVX1 U9644 ( .A(n17780), .Y(n16384) );
  INVX1 U9645 ( .A(n16387), .Y(n16385) );
  INVX1 U9646 ( .A(n16385), .Y(n16386) );
  AND2X1 U9647 ( .A(n17621), .B(n17615), .Y(n17501) );
  INVX1 U9648 ( .A(n17501), .Y(n16387) );
  INVX1 U9649 ( .A(n16390), .Y(n16388) );
  INVX1 U9650 ( .A(n16388), .Y(n16389) );
  BUFX2 U9651 ( .A(n18577), .Y(n16390) );
  INVX1 U9652 ( .A(n16393), .Y(n16391) );
  INVX1 U9653 ( .A(n16391), .Y(n16392) );
  AND2X1 U9654 ( .A(n16623), .B(n17114), .Y(n19768) );
  INVX1 U9655 ( .A(n19768), .Y(n16393) );
  INVX1 U9656 ( .A(n16396), .Y(n16394) );
  INVX1 U9657 ( .A(n16394), .Y(n16395) );
  BUFX2 U9658 ( .A(n18432), .Y(n16396) );
  INVX1 U9659 ( .A(n16399), .Y(n16397) );
  INVX1 U9660 ( .A(n16397), .Y(n16398) );
  AND2X2 U9661 ( .A(n17020), .B(n17627), .Y(n18359) );
  INVX1 U9662 ( .A(n18359), .Y(n16399) );
  INVX1 U9663 ( .A(n16402), .Y(n16400) );
  INVX1 U9664 ( .A(n16400), .Y(n16401) );
  BUFX2 U9665 ( .A(n18236), .Y(n16402) );
  INVX1 U9666 ( .A(n16405), .Y(n16403) );
  INVX1 U9667 ( .A(n16403), .Y(n16404) );
  AND2X1 U9668 ( .A(n17612), .B(n18175), .Y(n19767) );
  INVX1 U9669 ( .A(n19767), .Y(n16405) );
  INVX1 U9670 ( .A(n16408), .Y(n16406) );
  INVX1 U9671 ( .A(n16406), .Y(n16407) );
  AND2X1 U9672 ( .A(n18104), .B(n18405), .Y(n19774) );
  INVX1 U9673 ( .A(n19774), .Y(n16408) );
  INVX1 U9674 ( .A(n16411), .Y(n16409) );
  INVX1 U9675 ( .A(n16409), .Y(n16410) );
  AND2X2 U9676 ( .A(n19135), .B(n19134), .Y(n19167) );
  INVX1 U9677 ( .A(n19167), .Y(n16411) );
  INVX1 U9678 ( .A(n16414), .Y(n16412) );
  INVX1 U9679 ( .A(n16412), .Y(n16413) );
  AND2X1 U9680 ( .A(n18945), .B(n16416), .Y(n18783) );
  INVX1 U9681 ( .A(n18783), .Y(n16414) );
  INVX1 U9682 ( .A(n16417), .Y(n16415) );
  INVX1 U9683 ( .A(n16415), .Y(n16416) );
  AND2X1 U9684 ( .A(n18915), .B(n17078), .Y(n18806) );
  INVX1 U9685 ( .A(n18806), .Y(n16417) );
  INVX1 U9686 ( .A(n16420), .Y(n16418) );
  INVX1 U9687 ( .A(n16418), .Y(n16419) );
  AND2X1 U9688 ( .A(n17597), .B(n17467), .Y(n18297) );
  INVX1 U9689 ( .A(n18297), .Y(n16420) );
  INVX1 U9690 ( .A(n16423), .Y(n16421) );
  INVX1 U9691 ( .A(n16421), .Y(n16422) );
  AND2X1 U9692 ( .A(n19712), .B(n18155), .Y(n19771) );
  INVX1 U9693 ( .A(n19771), .Y(n16423) );
  INVX1 U9694 ( .A(n16426), .Y(n16424) );
  INVX1 U9695 ( .A(n16424), .Y(n16425) );
  AND2X2 U9696 ( .A(n18126), .B(n17013), .Y(n18148) );
  INVX1 U9697 ( .A(n18148), .Y(n16426) );
  INVX1 U9698 ( .A(n16429), .Y(n16427) );
  INVX1 U9699 ( .A(n16427), .Y(n16428) );
  BUFX2 U9700 ( .A(n19338), .Y(n16429) );
  INVX1 U9701 ( .A(n16432), .Y(n16430) );
  INVX1 U9702 ( .A(n16430), .Y(n16431) );
  OR2X1 U9703 ( .A(n17525), .B(n16521), .Y(n17553) );
  INVX1 U9704 ( .A(n17553), .Y(n16432) );
  INVX1 U9705 ( .A(n16435), .Y(n16433) );
  INVX1 U9706 ( .A(n16433), .Y(n16434) );
  AND2X1 U9707 ( .A(\lamb/scale_ts3/genblk1[2].mult/added[2] ), .B(n16571), 
        .Y(n19032) );
  INVX1 U9708 ( .A(n19032), .Y(n16435) );
  INVX1 U9709 ( .A(n16438), .Y(n16436) );
  INVX1 U9710 ( .A(n16436), .Y(n16437) );
  AND2X1 U9711 ( .A(n17759), .B(n17042), .Y(n17788) );
  INVX1 U9712 ( .A(n17788), .Y(n16438) );
  INVX1 U9713 ( .A(n16441), .Y(n16439) );
  INVX1 U9714 ( .A(n16439), .Y(n16440) );
  BUFX2 U9715 ( .A(n18515), .Y(n16441) );
  INVX1 U9716 ( .A(n16444), .Y(n16442) );
  INVX1 U9717 ( .A(n16442), .Y(n16443) );
  OR2X1 U9718 ( .A(\lamb/scale_ts0/genblk1[0].mult/added[3] ), .B(n17618), .Y(
        n17639) );
  INVX1 U9719 ( .A(n17639), .Y(n16444) );
  INVX1 U9720 ( .A(n16447), .Y(n16445) );
  INVX1 U9721 ( .A(n16445), .Y(n16446) );
  OR2X1 U9722 ( .A(\add_x_52/n1 ), .B(
        \lamb/scale_ls3/genblk1[1].mult/added[4] ), .Y(n18508) );
  INVX1 U9723 ( .A(n18508), .Y(n16447) );
  INVX1 U9724 ( .A(n16450), .Y(n16448) );
  INVX1 U9725 ( .A(n16448), .Y(n16449) );
  AND2X2 U9726 ( .A(n18763), .B(n16762), .Y(n18953) );
  INVX1 U9727 ( .A(n18953), .Y(n16450) );
  INVX1 U9728 ( .A(n16453), .Y(n16451) );
  INVX1 U9729 ( .A(n16451), .Y(n16452) );
  BUFX2 U9730 ( .A(n17486), .Y(n16453) );
  INVX1 U9731 ( .A(n16456), .Y(n16454) );
  INVX1 U9732 ( .A(n16454), .Y(n16455) );
  BUFX2 U9733 ( .A(n19289), .Y(n16456) );
  INVX1 U9734 ( .A(n16459), .Y(n16457) );
  INVX1 U9735 ( .A(n16457), .Y(n16458) );
  OR2X1 U9736 ( .A(\lamb/scale_ts1/genblk1[2].mult/added[4] ), .B(
        \add_x_68/n1 ), .Y(n17702) );
  INVX1 U9737 ( .A(n17702), .Y(n16459) );
  INVX1 U9738 ( .A(n16462), .Y(n16460) );
  INVX1 U9739 ( .A(n16460), .Y(n16461) );
  BUFX2 U9740 ( .A(n19333), .Y(n16462) );
  INVX1 U9741 ( .A(n16465), .Y(n16463) );
  INVX1 U9742 ( .A(n16463), .Y(n16464) );
  AND2X1 U9743 ( .A(n18348), .B(n19719), .Y(n19717) );
  INVX1 U9744 ( .A(n19717), .Y(n16465) );
  INVX1 U9745 ( .A(n16468), .Y(n16466) );
  INVX1 U9746 ( .A(n16466), .Y(n16467) );
  AND2X2 U9747 ( .A(n17036), .B(n17549), .Y(n17529) );
  INVX1 U9748 ( .A(n17529), .Y(n16468) );
  INVX1 U9749 ( .A(n16471), .Y(n16469) );
  INVX1 U9750 ( .A(n16469), .Y(n16470) );
  AND2X1 U9751 ( .A(n16554), .B(n16724), .Y(n18845) );
  INVX1 U9752 ( .A(n18845), .Y(n16471) );
  INVX1 U9753 ( .A(n16474), .Y(n16472) );
  INVX1 U9754 ( .A(n16472), .Y(n16473) );
  OR2X1 U9755 ( .A(n18898), .B(n17078), .Y(n18900) );
  INVX1 U9756 ( .A(n18900), .Y(n16474) );
  INVX1 U9757 ( .A(n16477), .Y(n16475) );
  INVX1 U9758 ( .A(n16475), .Y(n16476) );
  AND2X1 U9759 ( .A(\lamb/scale_ts1/genblk1[3].mult/added[3] ), .B(n17324), 
        .Y(n17327) );
  INVX1 U9760 ( .A(n17327), .Y(n16477) );
  INVX1 U9761 ( .A(n16480), .Y(n16478) );
  INVX1 U9762 ( .A(n16478), .Y(n16479) );
  AND2X1 U9763 ( .A(n18303), .B(n16576), .Y(n18289) );
  INVX1 U9764 ( .A(n18289), .Y(n16480) );
  INVX1 U9765 ( .A(n16483), .Y(n16481) );
  INVX1 U9766 ( .A(n16481), .Y(n16482) );
  AND2X1 U9767 ( .A(n18323), .B(n18322), .Y(n18331) );
  INVX1 U9768 ( .A(n18331), .Y(n16483) );
  INVX1 U9769 ( .A(n16486), .Y(n16484) );
  INVX1 U9770 ( .A(n16484), .Y(n16485) );
  AND2X1 U9771 ( .A(n17594), .B(n17589), .Y(n17391) );
  INVX1 U9772 ( .A(n17391), .Y(n16486) );
  INVX1 U9773 ( .A(n16489), .Y(n16487) );
  INVX1 U9774 ( .A(n16487), .Y(n16488) );
  AND2X1 U9775 ( .A(n17616), .B(n16611), .Y(n17648) );
  INVX1 U9776 ( .A(n17648), .Y(n16489) );
  INVX1 U9777 ( .A(n16492), .Y(n16490) );
  INVX1 U9778 ( .A(n16490), .Y(n16491) );
  AND2X1 U9779 ( .A(\lamb/scale_ls2/genblk1[1].mult/added[2] ), .B(
        \lamb/scale_ls2/genblk1[1].mult/added[1] ), .Y(n18151) );
  INVX1 U9780 ( .A(n18151), .Y(n16492) );
  INVX1 U9781 ( .A(n16495), .Y(n16493) );
  INVX1 U9782 ( .A(n16493), .Y(n16494) );
  AND2X1 U9783 ( .A(n19219), .B(n19220), .Y(n19242) );
  INVX1 U9784 ( .A(n19242), .Y(n16495) );
  INVX1 U9785 ( .A(n16498), .Y(n16496) );
  INVX1 U9786 ( .A(n16496), .Y(n16497) );
  OR2X1 U9787 ( .A(n16734), .B(n19726), .Y(n19659) );
  INVX1 U9788 ( .A(n19659), .Y(n16498) );
  INVX1 U9789 ( .A(n16501), .Y(n16499) );
  INVX1 U9790 ( .A(n16499), .Y(n16500) );
  AND2X1 U9791 ( .A(n19246), .B(n16527), .Y(n19511) );
  INVX1 U9792 ( .A(n19511), .Y(n16501) );
  INVX1 U9793 ( .A(n16504), .Y(n16502) );
  INVX1 U9794 ( .A(n16502), .Y(n16503) );
  OR2X1 U9795 ( .A(n17759), .B(n16629), .Y(n17792) );
  INVX1 U9796 ( .A(n17792), .Y(n16504) );
  INVX1 U9797 ( .A(n16507), .Y(n16505) );
  INVX1 U9798 ( .A(n16505), .Y(n16506) );
  AND2X2 U9799 ( .A(n19256), .B(n18776), .Y(n18787) );
  INVX1 U9800 ( .A(n18787), .Y(n16507) );
  INVX1 U9801 ( .A(n16510), .Y(n16508) );
  INVX1 U9802 ( .A(n16508), .Y(n16509) );
  AND2X1 U9803 ( .A(\lamb/scale_ts1/genblk1[2].mult/added[4] ), .B(
        \add_x_68/n1 ), .Y(n17659) );
  INVX1 U9804 ( .A(n17659), .Y(n16510) );
  INVX1 U9805 ( .A(n16513), .Y(n16511) );
  INVX1 U9806 ( .A(n16511), .Y(n16512) );
  AND2X1 U9807 ( .A(n18915), .B(n18945), .Y(n18916) );
  INVX1 U9808 ( .A(n18916), .Y(n16513) );
  INVX1 U9809 ( .A(n16516), .Y(n16514) );
  INVX1 U9810 ( .A(n16514), .Y(n16515) );
  OR2X2 U9811 ( .A(n18427), .B(n18426), .Y(n18444) );
  INVX1 U9812 ( .A(n18444), .Y(n16516) );
  INVX1 U9813 ( .A(n16519), .Y(n16517) );
  INVX1 U9814 ( .A(n16517), .Y(n16518) );
  INVX1 U9815 ( .A(n17700), .Y(n16519) );
  INVX1 U9816 ( .A(n16522), .Y(n16520) );
  INVX1 U9817 ( .A(n16520), .Y(n16521) );
  BUFX2 U9818 ( .A(n17521), .Y(n16522) );
  INVX1 U9819 ( .A(n16525), .Y(n16523) );
  INVX1 U9820 ( .A(n16523), .Y(n16524) );
  OR2X1 U9821 ( .A(\lamb/scale_ts0/genblk1[1].mult/added[3] ), .B(n16934), .Y(
        n17425) );
  INVX1 U9822 ( .A(n17425), .Y(n16525) );
  INVX1 U9823 ( .A(n16528), .Y(n16526) );
  INVX1 U9824 ( .A(n16526), .Y(n16527) );
  BUFX2 U9825 ( .A(n19251), .Y(n16528) );
  INVX1 U9826 ( .A(n16531), .Y(n16529) );
  INVX1 U9827 ( .A(n16529), .Y(n16530) );
  BUFX2 U9828 ( .A(n17880), .Y(n16531) );
  INVX1 U9829 ( .A(n16534), .Y(n16532) );
  INVX1 U9830 ( .A(n16532), .Y(n16533) );
  BUFX2 U9831 ( .A(n18584), .Y(n16534) );
  INVX1 U9832 ( .A(n16537), .Y(n16535) );
  INVX1 U9833 ( .A(n16535), .Y(n16536) );
  BUFX2 U9834 ( .A(n19534), .Y(n16537) );
  INVX1 U9835 ( .A(n16540), .Y(n16538) );
  INVX1 U9836 ( .A(n16538), .Y(n16539) );
  BUFX2 U9837 ( .A(n19537), .Y(n16540) );
  INVX1 U9838 ( .A(n16543), .Y(n16541) );
  INVX1 U9839 ( .A(n16541), .Y(n16542) );
  BUFX2 U9840 ( .A(n19540), .Y(n16543) );
  INVX1 U9841 ( .A(n16546), .Y(n16544) );
  INVX1 U9842 ( .A(n16544), .Y(n16545) );
  BUFX2 U9843 ( .A(n19542), .Y(n16546) );
  INVX1 U9844 ( .A(n16549), .Y(n16547) );
  INVX1 U9845 ( .A(n16547), .Y(n16548) );
  AND2X1 U9846 ( .A(n17222), .B(n17588), .Y(n17369) );
  INVX1 U9847 ( .A(n17369), .Y(n16549) );
  INVX1 U9848 ( .A(n16552), .Y(n16550) );
  INVX1 U9849 ( .A(n16550), .Y(n16551) );
  AND2X1 U9850 ( .A(n18821), .B(n18822), .Y(n18828) );
  INVX1 U9851 ( .A(n18828), .Y(n16552) );
  INVX1 U9852 ( .A(n16555), .Y(n16553) );
  INVX1 U9853 ( .A(n16553), .Y(n16554) );
  BUFX2 U9854 ( .A(n18859), .Y(n16555) );
  INVX1 U9855 ( .A(n16556), .Y(n18859) );
  INVX1 U9856 ( .A(n18817), .Y(n16557) );
  INVX1 U9857 ( .A(n18957), .Y(n16558) );
  INVX1 U9858 ( .A(n18818), .Y(n16559) );
  NOR2X1 U9859 ( .A(n16559), .B(n16560), .Y(n16556) );
  NOR2X1 U9860 ( .A(n16557), .B(n16558), .Y(n16561) );
  INVX1 U9861 ( .A(n16561), .Y(n16560) );
  INVX1 U9862 ( .A(n16564), .Y(n16562) );
  INVX1 U9863 ( .A(n16562), .Y(n16563) );
  AND2X2 U9864 ( .A(n16763), .B(n18763), .Y(n18795) );
  INVX1 U9865 ( .A(n18795), .Y(n16564) );
  INVX1 U9866 ( .A(n16567), .Y(n16565) );
  INVX1 U9867 ( .A(n16565), .Y(n16566) );
  BUFX2 U9868 ( .A(n18501), .Y(n16567) );
  OR2X1 U9869 ( .A(n17095), .B(\lamb/scale_ts0/genblk1[2].mult/added[2] ), .Y(
        n17265) );
  AND2X1 U9870 ( .A(n18752), .B(n17028), .Y(
        \lamb/scale_ts1/genblk1[0].mult/logA[1] ) );
  AND2X1 U9871 ( .A(n16645), .B(n18287), .Y(n18270) );
  XOR2X1 U9872 ( .A(n17594), .B(n16859), .Y(n18322) );
  OR2X1 U9873 ( .A(n17045), .B(n17966), .Y(n17985) );
  AND2X1 U9874 ( .A(n16629), .B(n17759), .Y(n17777) );
  AND2X1 U9875 ( .A(n17124), .B(n17628), .Y(
        \lamb/scale_bs2/genblk1[0].mult/logA[2] ) );
  AND2X1 U9876 ( .A(n18303), .B(n17068), .Y(
        \lamb/scale_ls2/genblk1[0].mult/logA[1] ) );
  AND2X1 U9877 ( .A(n16745), .B(n19726), .Y(n18294) );
  AND2X1 U9878 ( .A(n17062), .B(n17029), .Y(n18243) );
  AND2X1 U9879 ( .A(n16896), .B(n16980), .Y(n19742) );
  AND2X1 U9880 ( .A(n19666), .B(n16578), .Y(n17362) );
  OR2X1 U9881 ( .A(n16757), .B(n16655), .Y(n17847) );
  OR2X1 U9882 ( .A(n19267), .B(n16981), .Y(n19273) );
  AND2X1 U9883 ( .A(n18414), .B(n17031), .Y(
        \lamb/scale_bs3/genblk1[0].mult/logA[3] ) );
  AND2X1 U9884 ( .A(n17004), .B(n18171), .Y(n18173) );
  AND2X1 U9885 ( .A(n16642), .B(n16891), .Y(n17580) );
  AND2X1 U9886 ( .A(n18414), .B(n17124), .Y(n9909) );
  OR2X1 U9887 ( .A(n17741), .B(n16590), .Y(n17755) );
  AND2X1 U9888 ( .A(n19332), .B(n16624), .Y(n19334) );
  OR2X1 U9889 ( .A(n19274), .B(n17043), .Y(n19277) );
  AND2X1 U9890 ( .A(n17068), .B(n17630), .Y(
        \lamb/scale_ts1/genblk1[3].mult/logA[1] ) );
  OR2X1 U9891 ( .A(n16901), .B(n18526), .Y(n18524) );
  AND2X1 U9892 ( .A(n16637), .B(n17055), .Y(n19072) );
  AND2X1 U9893 ( .A(n16995), .B(n16643), .Y(n19266) );
  OR2X1 U9894 ( .A(n16806), .B(n18435), .Y(n18497) );
  AND2X1 U9895 ( .A(n18434), .B(n16639), .Y(n18436) );
  AND2X1 U9896 ( .A(n17094), .B(n17749), .Y(n17743) );
  OR2X1 U9897 ( .A(n17055), .B(n19053), .Y(n19040) );
  OR2X1 U9898 ( .A(n19193), .B(n17083), .Y(n19166) );
  OR2X1 U9899 ( .A(n19148), .B(n17027), .Y(n19149) );
  AND2X1 U9900 ( .A(n18882), .B(n16641), .Y(n18875) );
  AND2X1 U9901 ( .A(n16748), .B(n16735), .Y(n18897) );
  OR2X1 U9902 ( .A(n18938), .B(n17073), .Y(n18917) );
  AND2X1 U9903 ( .A(n18929), .B(n16930), .Y(n19548) );
  AND2X1 U9904 ( .A(n16626), .B(n18757), .Y(n18769) );
  OR2X1 U9905 ( .A(n16620), .B(n17101), .Y(n19544) );
  OR2X1 U9906 ( .A(n17096), .B(n16569), .Y(n19543) );
  OR2X1 U9907 ( .A(n16568), .B(n16703), .Y(n19566) );
  OR2X1 U9908 ( .A(n16569), .B(n16703), .Y(n19588) );
  OR2X1 U9909 ( .A(n16569), .B(n16704), .Y(n19653) );
  OR2X1 U9910 ( .A(n16568), .B(n16704), .Y(n19616) );
  OR2X1 U9911 ( .A(n17096), .B(n16568), .Y(n19520) );
  AND2X1 U9912 ( .A(n16572), .B(n18070), .Y(n18081) );
  AND2X1 U9913 ( .A(n16632), .B(n18018), .Y(n19705) );
  AND2X1 U9914 ( .A(n16758), .B(n16747), .Y(n17836) );
  AND2X1 U9915 ( .A(n16752), .B(n19620), .Y(n19606) );
  INVX1 U9916 ( .A(n19606), .Y(n16568) );
  AND2X1 U9917 ( .A(n19620), .B(n16751), .Y(n19639) );
  INVX1 U9918 ( .A(n19639), .Y(n16569) );
  AND2X1 U9919 ( .A(n17578), .B(n17579), .Y(n17584) );
  INVX1 U9920 ( .A(n17584), .Y(n16570) );
  AND2X1 U9921 ( .A(n18963), .B(n18962), .Y(n19005) );
  INVX1 U9922 ( .A(n19005), .Y(n16571) );
  AND2X1 U9923 ( .A(\lamb/scale_ts2/genblk1[3].mult/added[3] ), .B(n18082), 
        .Y(n18069) );
  INVX1 U9924 ( .A(n18069), .Y(n16572) );
  BUFX2 U9925 ( .A(n18092), .Y(n16573) );
  AND2X1 U9926 ( .A(n18234), .B(n18226), .Y(n18227) );
  INVX1 U9927 ( .A(n18227), .Y(n16574) );
  AND2X1 U9928 ( .A(n19210), .B(n19214), .Y(n19236) );
  INVX1 U9929 ( .A(n19236), .Y(n16575) );
  BUFX2 U9930 ( .A(n18749), .Y(n16576) );
  AND2X1 U9931 ( .A(n19262), .B(n19283), .Y(n19310) );
  INVX1 U9932 ( .A(n19310), .Y(n16577) );
  OR2X1 U9933 ( .A(n18337), .B(n18334), .Y(n19667) );
  INVX1 U9934 ( .A(n19667), .Y(n16578) );
  AND2X1 U9935 ( .A(n18937), .B(n19547), .Y(n19623) );
  INVX1 U9936 ( .A(n19623), .Y(n16579) );
  AND2X1 U9937 ( .A(n18937), .B(n16512), .Y(n19570) );
  INVX1 U9938 ( .A(n19570), .Y(n16580) );
  AND2X1 U9939 ( .A(n19073), .B(n16637), .Y(n19054) );
  INVX1 U9940 ( .A(n19054), .Y(n16581) );
  BUFX2 U9941 ( .A(n17357), .Y(n16582) );
  OR2X1 U9942 ( .A(n16763), .B(n18905), .Y(n19269) );
  INVX1 U9943 ( .A(n19269), .Y(n16583) );
  AND2X1 U9944 ( .A(n16660), .B(n18923), .Y(n18937) );
  INVX1 U9945 ( .A(n18937), .Y(n16584) );
  OR2X1 U9946 ( .A(n16395), .B(n16926), .Y(n18551) );
  INVX1 U9947 ( .A(n18551), .Y(n16585) );
  BUFX2 U9948 ( .A(n17677), .Y(n16586) );
  AND2X1 U9949 ( .A(n17046), .B(n16554), .Y(n18836) );
  INVX1 U9950 ( .A(n18836), .Y(n16587) );
  BUFX2 U9951 ( .A(n18113), .Y(n16588) );
  BUFX2 U9952 ( .A(n17869), .Y(n16589) );
  BUFX2 U9953 ( .A(n17742), .Y(n16590) );
  BUFX2 U9954 ( .A(n17398), .Y(n16591) );
  BUFX2 U9955 ( .A(n17191), .Y(n16592) );
  BUFX2 U9956 ( .A(n17193), .Y(n16593) );
  BUFX2 U9957 ( .A(n19247), .Y(n16594) );
  BUFX2 U9958 ( .A(n19231), .Y(n16595) );
  BUFX2 U9959 ( .A(n19672), .Y(n16596) );
  AND2X1 U9960 ( .A(n18413), .B(n19693), .Y(n19694) );
  INVX1 U9961 ( .A(n19694), .Y(n16597) );
  AND2X1 U9962 ( .A(n18020), .B(n18018), .Y(n19706) );
  INVX1 U9963 ( .A(n19706), .Y(n16598) );
  INVX1 U9964 ( .A(n17747), .Y(n16599) );
  AND2X1 U9965 ( .A(n17961), .B(n18003), .Y(n18007) );
  INVX1 U9966 ( .A(n18007), .Y(n16600) );
  AND2X1 U9967 ( .A(n16750), .B(n18217), .Y(n18223) );
  INVX1 U9968 ( .A(n18223), .Y(n16601) );
  AND2X1 U9969 ( .A(n19099), .B(n19134), .Y(n19192) );
  INVX1 U9970 ( .A(n19192), .Y(n16602) );
  BUFX2 U9971 ( .A(n17492), .Y(n16603) );
  AND2X1 U9972 ( .A(n19053), .B(n19052), .Y(n19071) );
  INVX1 U9973 ( .A(n19071), .Y(n16604) );
  AND2X1 U9974 ( .A(n17499), .B(n17498), .Y(n17504) );
  INVX1 U9975 ( .A(n17504), .Y(n16605) );
  BUFX2 U9976 ( .A(n19190), .Y(n16606) );
  AND2X1 U9977 ( .A(n19210), .B(n19209), .Y(n19234) );
  INVX1 U9978 ( .A(n19234), .Y(n16607) );
  BUFX2 U9979 ( .A(n18149), .Y(n16608) );
  AND2X1 U9980 ( .A(n16452), .B(n17485), .Y(n17494) );
  INVX1 U9981 ( .A(n17494), .Y(n16609) );
  OR2X1 U9982 ( .A(n18186), .B(n18434), .Y(n18193) );
  INVX1 U9983 ( .A(n18193), .Y(n16610) );
  AND2X1 U9984 ( .A(\lamb/scale_ts0/genblk1[0].mult/added[3] ), .B(n17623), 
        .Y(n17635) );
  INVX1 U9985 ( .A(n17635), .Y(n16611) );
  OR2X1 U9986 ( .A(n16618), .B(n19267), .Y(n19265) );
  INVX1 U9987 ( .A(n19265), .Y(n16612) );
  BUFX2 U9988 ( .A(n17490), .Y(n16613) );
  OR2X1 U9989 ( .A(n16542), .B(n17051), .Y(n19613) );
  INVX1 U9990 ( .A(n19613), .Y(n16614) );
  OR2X1 U9991 ( .A(n19225), .B(n19230), .Y(n19240) );
  INVX1 U9992 ( .A(n19240), .Y(n16615) );
  OR2X1 U9993 ( .A(n16545), .B(n17051), .Y(n19617) );
  INVX1 U9994 ( .A(n19617), .Y(n16616) );
  BUFX2 U9995 ( .A(n18181), .Y(n16617) );
  OR2X1 U9996 ( .A(n16551), .B(n18823), .Y(n19262) );
  INVX1 U9997 ( .A(n19262), .Y(n16618) );
  AND2X1 U9998 ( .A(n17609), .B(n19703), .Y(n17948) );
  INVX1 U9999 ( .A(n17948), .Y(n16619) );
  AND2X1 U10000 ( .A(n18754), .B(n18906), .Y(n19256) );
  INVX1 U10001 ( .A(n19256), .Y(n16620) );
  AND2X1 U10002 ( .A(n19310), .B(n19286), .Y(n19313) );
  INVX1 U10003 ( .A(n19313), .Y(n16621) );
  AND2X1 U10004 ( .A(n17598), .B(n17602), .Y(n17585) );
  INVX1 U10005 ( .A(n17585), .Y(n16622) );
  BUFX2 U10006 ( .A(n18180), .Y(n16623) );
  AND2X1 U10007 ( .A(n17101), .B(n19329), .Y(n19335) );
  INVX1 U10008 ( .A(n19335), .Y(n16624) );
  AND2X1 U10009 ( .A(n16626), .B(n18791), .Y(n18943) );
  INVX1 U10010 ( .A(n18943), .Y(n16625) );
  AND2X1 U10011 ( .A(n18734), .B(n18733), .Y(n18784) );
  INVX1 U10012 ( .A(n18784), .Y(n16626) );
  BUFX2 U10013 ( .A(n17645), .Y(n16627) );
  AND2X1 U10014 ( .A(\lamb/scale_ts1/genblk1[0].mult/added[2] ), .B(
        \lamb/scale_ts1/genblk1[0].mult/added[1] ), .Y(n17489) );
  INVX1 U10015 ( .A(n17489), .Y(n16628) );
  OR2X1 U10016 ( .A(\lamb/scale_ds1/genblk1[1].mult/added[4] ), .B(
        \add_x_73/n1 ), .Y(n17827) );
  INVX1 U10017 ( .A(n17827), .Y(n16629) );
  AND2X1 U10018 ( .A(\lamb/scale_ds2/genblk1[3].mult/added[1] ), .B(
        \lamb/scale_ds2/genblk1[3].mult/added[2] ), .Y(n18091) );
  INVX1 U10019 ( .A(n18091), .Y(n16630) );
  OR2X1 U10020 ( .A(n16629), .B(n16437), .Y(n17825) );
  INVX1 U10021 ( .A(n17825), .Y(n16631) );
  BUFX2 U10022 ( .A(n18019), .Y(n16632) );
  OR2X1 U10023 ( .A(n16536), .B(n17051), .Y(n19607) );
  INVX1 U10024 ( .A(n19607), .Y(n16633) );
  OR2X1 U10025 ( .A(n16539), .B(n17051), .Y(n19610) );
  INVX1 U10026 ( .A(n19610), .Y(n16634) );
  AND2X1 U10027 ( .A(n19215), .B(n19204), .Y(n19235) );
  INVX1 U10028 ( .A(n19235), .Y(n16635) );
  BUFX2 U10029 ( .A(n17542), .Y(n16636) );
  AND2X1 U10030 ( .A(n19058), .B(n19061), .Y(n19070) );
  INVX1 U10031 ( .A(n19070), .Y(n16637) );
  AND2X1 U10032 ( .A(n17630), .B(n16921), .Y(n17451) );
  INVX1 U10033 ( .A(n17451), .Y(n16638) );
  AND2X1 U10034 ( .A(n16647), .B(n18190), .Y(n18433) );
  INVX1 U10035 ( .A(n18433), .Y(n16639) );
  INVX1 U10036 ( .A(n18531), .Y(n16640) );
  AND2X1 U10037 ( .A(n18850), .B(n18849), .Y(n18867) );
  INVX1 U10038 ( .A(n18867), .Y(n16641) );
  AND2X1 U10039 ( .A(n17578), .B(n17222), .Y(n17582) );
  INVX1 U10040 ( .A(n17582), .Y(n16642) );
  AND2X1 U10041 ( .A(n19264), .B(n19270), .Y(n19280) );
  INVX1 U10042 ( .A(n19280), .Y(n16643) );
  AND2X1 U10043 ( .A(n19264), .B(n18766), .Y(n18788) );
  INVX1 U10044 ( .A(n18788), .Y(n16644) );
  OR2X1 U10045 ( .A(n18268), .B(n17495), .Y(n18283) );
  INVX1 U10046 ( .A(n18283), .Y(n16645) );
  BUFX2 U10047 ( .A(n17900), .Y(n16646) );
  BUFX2 U10048 ( .A(n18183), .Y(n16647) );
  BUFX2 U10049 ( .A(n19282), .Y(n16648) );
  BUFX2 U10050 ( .A(n18008), .Y(n16649) );
  OR2X1 U10051 ( .A(n16750), .B(n16760), .Y(n18218) );
  INVX1 U10052 ( .A(n18218), .Y(n16650) );
  AND2X1 U10053 ( .A(n18911), .B(n18910), .Y(n19342) );
  INVX1 U10054 ( .A(n19342), .Y(n16651) );
  BUFX2 U10055 ( .A(n17444), .Y(n16652) );
  AND2X1 U10056 ( .A(n18309), .B(n17665), .Y(n19754) );
  INVX1 U10057 ( .A(n19754), .Y(n16653) );
  BUFX2 U10058 ( .A(n17801), .Y(n16654) );
  BUFX2 U10059 ( .A(n17842), .Y(n16655) );
  BUFX2 U10060 ( .A(n19129), .Y(n16656) );
  AND2X1 U10061 ( .A(n19264), .B(n16449), .Y(n19257) );
  INVX1 U10062 ( .A(n19257), .Y(n16657) );
  AND2X1 U10063 ( .A(n18938), .B(n17073), .Y(n18945) );
  INVX1 U10064 ( .A(n18945), .Y(n16658) );
  BUFX2 U10065 ( .A(n17311), .Y(n16659) );
  OR2X1 U10066 ( .A(n17107), .B(n18905), .Y(n18921) );
  INVX1 U10067 ( .A(n18921), .Y(n16660) );
  AND2X1 U10068 ( .A(n18752), .B(n16419), .Y(n18303) );
  INVX1 U10069 ( .A(n18303), .Y(n16661) );
  BUFX2 U10070 ( .A(n19028), .Y(n16662) );
  BUFX2 U10071 ( .A(n18212), .Y(n16663) );
  AND2X1 U10072 ( .A(n17597), .B(n17630), .Y(n17738) );
  INVX1 U10073 ( .A(n17738), .Y(n16664) );
  BUFX2 U10074 ( .A(n18580), .Y(n16665) );
  BUFX2 U10075 ( .A(n19064), .Y(n16666) );
  BUFX2 U10076 ( .A(n17135), .Y(n16667) );
  BUFX2 U10077 ( .A(n17151), .Y(n16668) );
  BUFX2 U10078 ( .A(n17157), .Y(n16669) );
  BUFX2 U10079 ( .A(\lamb/scale_ls3/genblk1[1].mult/logA[2] ), .Y(n16670) );
  BUFX2 U10080 ( .A(\lamb/scale_ts1/genblk1[1].mult/logA[1] ), .Y(n16671) );
  BUFX2 U10081 ( .A(\lamb/scale_ds1/genblk1[1].mult/logA[1] ), .Y(n16672) );
  BUFX2 U10082 ( .A(\lamb/scale_ts0/genblk1[1].mult/logA[2] ), .Y(n16673) );
  BUFX2 U10083 ( .A(n19345), .Y(n16674) );
  BUFX2 U10084 ( .A(n19430), .Y(n16675) );
  BUFX2 U10085 ( .A(n19673), .Y(n16676) );
  BUFX2 U10086 ( .A(\lamb/scale_ts2/genblk1[1].mult/logA[1] ), .Y(n16677) );
  BUFX2 U10087 ( .A(\lamb/scale_ts3/genblk1[3].mult/logA[2] ), .Y(n16678) );
  BUFX2 U10088 ( .A(\lamb/scale_ds3/genblk1[3].mult/logA[2] ), .Y(n16679) );
  BUFX2 U10089 ( .A(\lamb/scale_ds3/genblk1[2].mult/logA[1] ), .Y(n16680) );
  BUFX2 U10090 ( .A(\lamb/scale_ds3/genblk1[2].mult/logA[2] ), .Y(n16681) );
  BUFX2 U10091 ( .A(\lamb/scale_ls3/genblk1[2].mult/logA[0] ), .Y(n16682) );
  BUFX2 U10092 ( .A(\lamb/scale_ls3/genblk1[1].mult/logA[1] ), .Y(n16683) );
  BUFX2 U10093 ( .A(\lamb/scale_ls3/genblk1[0].mult/logA[1] ), .Y(n16684) );
  BUFX2 U10094 ( .A(\lamb/scale_ls3/genblk1[0].mult/logA[2] ), .Y(n16685) );
  BUFX2 U10095 ( .A(\lamb/scale_ts2/genblk1[3].mult/logA[1] ), .Y(n16686) );
  BUFX2 U10096 ( .A(\lamb/scale_ts2/genblk1[2].mult/logA[1] ), .Y(n16687) );
  OR2X1 U10097 ( .A(n17950), .B(n17949), .Y(n17653) );
  BUFX2 U10098 ( .A(\lamb/scale_ts2/genblk1[1].mult/logA[2] ), .Y(n16688) );
  BUFX2 U10099 ( .A(\lamb/scale_ds2/genblk1[3].mult/logA[1] ), .Y(n16689) );
  BUFX2 U10100 ( .A(\lamb/scale_ds2/genblk1[2].mult/logA[1] ), .Y(n16690) );
  BUFX2 U10101 ( .A(\lamb/scale_ds2/genblk1[2].mult/logA[2] ), .Y(n16691) );
  BUFX2 U10102 ( .A(\lamb/scale_ds2/genblk1[1].mult/logA[1] ), .Y(n16692) );
  BUFX2 U10103 ( .A(\lamb/scale_ls2/genblk1[0].mult/logA[2] ), .Y(n16693) );
  BUFX2 U10104 ( .A(\lamb/scale_ts1/genblk1[2].mult/logA[2] ), .Y(n16694) );
  BUFX2 U10105 ( .A(\lamb/scale_ts0/genblk1[1].mult/logA[1] ), .Y(n16695) );
  BUFX2 U10106 ( .A(n19076), .Y(n16696) );
  BUFX2 U10107 ( .A(n19248), .Y(n16697) );
  BUFX2 U10108 ( .A(n16304), .Y(n16698) );
  INVX1 U10109 ( .A(n16311), .Y(n16699) );
  AND2X1 U10110 ( .A(n19737), .B(n19736), .Y(n16311) );
  INVX1 U10111 ( .A(n16309), .Y(n16700) );
  OR2X1 U10112 ( .A(n19748), .B(n19747), .Y(n16309) );
  INVX1 U10113 ( .A(n16308), .Y(n16701) );
  OR2X1 U10114 ( .A(n19750), .B(n19749), .Y(n16308) );
  INVX1 U10115 ( .A(n18366), .Y(n16702) );
  AND2X1 U10116 ( .A(n18369), .B(n16886), .Y(n18366) );
  INVX1 U10117 ( .A(n19581), .Y(n16703) );
  AND2X1 U10118 ( .A(n17096), .B(n19591), .Y(n19581) );
  INVX1 U10119 ( .A(n19638), .Y(n16704) );
  AND2X1 U10120 ( .A(n19593), .B(n17096), .Y(n19638) );
  INVX1 U10121 ( .A(n19531), .Y(n16705) );
  OR2X1 U10122 ( .A(n16762), .B(n19523), .Y(n19531) );
  INVX1 U10123 ( .A(n19635), .Y(n16706) );
  OR2X1 U10124 ( .A(n16579), .B(n19622), .Y(n19635) );
  INVX1 U10125 ( .A(n19520), .Y(n16707) );
  INVX1 U10126 ( .A(n19392), .Y(n16708) );
  OR2X1 U10127 ( .A(n19358), .B(n19356), .Y(n19392) );
  INVX1 U10128 ( .A(n16306), .Y(n16709) );
  OR2X1 U10129 ( .A(n16904), .B(n18298), .Y(n16306) );
  BUFX2 U10130 ( .A(\lamb/scale_ts0/genblk1[0].mult/logA[2] ), .Y(n16710) );
  BUFX2 U10131 ( .A(n17158), .Y(n16711) );
  BUFX2 U10132 ( .A(n17415), .Y(n16712) );
  INVX1 U10133 ( .A(n19068), .Y(n16713) );
  OR2X1 U10134 ( .A(n19063), .B(n19045), .Y(n19068) );
  BUFX2 U10135 ( .A(n17284), .Y(n16714) );
  INVX1 U10136 ( .A(n19077), .Y(n16715) );
  OR2X1 U10137 ( .A(n19042), .B(n16461), .Y(n19077) );
  BUFX2 U10138 ( .A(n17373), .Y(n16716) );
  BUFX2 U10139 ( .A(n19349), .Y(n16717) );
  INVX1 U10140 ( .A(n19616), .Y(n16718) );
  INVX1 U10141 ( .A(n19543), .Y(n16719) );
  INVX1 U10142 ( .A(n19566), .Y(n16720) );
  INVX1 U10143 ( .A(n19588), .Y(n16721) );
  INVX1 U10144 ( .A(n19653), .Y(n16722) );
  INVX1 U10145 ( .A(n18932), .Y(n16723) );
  AND2X1 U10146 ( .A(n18764), .B(n17073), .Y(n18932) );
  INVX1 U10147 ( .A(n16725), .Y(n16724) );
  INVX1 U10148 ( .A(n18798), .Y(n16726) );
  INVX1 U10149 ( .A(n18799), .Y(n16727) );
  INVX1 U10150 ( .A(n18800), .Y(n16728) );
  NOR2X1 U10151 ( .A(n16728), .B(n16729), .Y(n16725) );
  NOR2X1 U10152 ( .A(n16726), .B(n16727), .Y(n16730) );
  INVX1 U10153 ( .A(n16730), .Y(n16729) );
  INVX1 U10154 ( .A(n16732), .Y(n16731) );
  BUFX2 U10155 ( .A(n18235), .Y(n16732) );
  INVX1 U10156 ( .A(n16734), .Y(n16733) );
  BUFX2 U10157 ( .A(n19731), .Y(n16734) );
  INVX1 U10158 ( .A(n18944), .Y(n16735) );
  AND2X1 U10159 ( .A(n18945), .B(n18940), .Y(n18944) );
  INVX1 U10160 ( .A(n16737), .Y(n16736) );
  BUFX2 U10161 ( .A(n19595), .Y(n16737) );
  NAND2X1 U10162 ( .A(n16738), .B(n16739), .Y(n19595) );
  INVX1 U10163 ( .A(n16413), .Y(n16740) );
  NAND2X1 U10164 ( .A(n18788), .B(n17107), .Y(n16738) );
  NAND2X1 U10165 ( .A(n18788), .B(n16740), .Y(n16739) );
  BUFX2 U10166 ( .A(n17570), .Y(n16741) );
  INVX1 U10167 ( .A(n16743), .Y(n16742) );
  BUFX2 U10168 ( .A(n17839), .Y(n16743) );
  INVX1 U10169 ( .A(n16745), .Y(n16744) );
  BUFX2 U10170 ( .A(n19727), .Y(n16745) );
  INVX1 U10171 ( .A(n18413), .Y(n16746) );
  AND2X1 U10172 ( .A(n17630), .B(n16338), .Y(n18413) );
  BUFX2 U10173 ( .A(n17843), .Y(n16747) );
  BUFX2 U10174 ( .A(n18815), .Y(n16748) );
  INVX1 U10175 ( .A(n17912), .Y(n16749) );
  OR2X1 U10176 ( .A(\lamb/scale_ts2/genblk1[2].mult/added[4] ), .B(
        \add_x_55/n1 ), .Y(n17912) );
  BUFX2 U10177 ( .A(n18216), .Y(n16750) );
  INVX1 U10178 ( .A(n16752), .Y(n16751) );
  BUFX2 U10179 ( .A(n19621), .Y(n16752) );
  NOR2X1 U10180 ( .A(n16753), .B(n16754), .Y(n19621) );
  INVX1 U10181 ( .A(n18761), .Y(n16755) );
  INVX1 U10182 ( .A(n18762), .Y(n16756) );
  NOR2X1 U10183 ( .A(n16755), .B(n16756), .Y(n16753) );
  NOR2X1 U10184 ( .A(n19256), .B(n16736), .Y(n16754) );
  INVX1 U10185 ( .A(n16758), .Y(n16757) );
  BUFX2 U10186 ( .A(n17835), .Y(n16758) );
  INVX1 U10187 ( .A(n16760), .Y(n16759) );
  BUFX2 U10188 ( .A(n18222), .Y(n16760) );
  BUFX2 U10189 ( .A(n18224), .Y(n16761) );
  INVX1 U10190 ( .A(n16763), .Y(n16762) );
  BUFX2 U10191 ( .A(n18954), .Y(n16763) );
  INVX1 U10192 ( .A(n16765), .Y(n16764) );
  INVX1 U10193 ( .A(n16361), .Y(n16766) );
  INVX1 U10194 ( .A(n18590), .Y(n16767) );
  NOR2X1 U10195 ( .A(n16767), .B(n16768), .Y(n16765) );
  NOR2X1 U10196 ( .A(n18588), .B(n16766), .Y(n16769) );
  INVX1 U10197 ( .A(n16769), .Y(n16768) );
  BUFX2 U10198 ( .A(n9917), .Y(n16770) );
  NOR2X1 U10199 ( .A(n16771), .B(n16772), .Y(n9917) );
  INVX1 U10200 ( .A(n16497), .Y(n16773) );
  NOR2X1 U10201 ( .A(n17120), .B(n16773), .Y(n16771) );
  INVX1 U10202 ( .A(n19657), .Y(n16774) );
  INVX1 U10203 ( .A(n19658), .Y(n16775) );
  NOR2X1 U10204 ( .A(n16774), .B(n16775), .Y(n16772) );
  BUFX2 U10205 ( .A(\lamb/scale_ts1/genblk1[0].mult/logB[1] ), .Y(n16776) );
  BUFX2 U10206 ( .A(\lamb/scale_ls3/genblk1[0].mult/logB[1] ), .Y(n16777) );
  NOR2X1 U10207 ( .A(n16778), .B(n16779), .Y(
        \lamb/scale_ls3/genblk1[0].mult/logB[1] ) );
  NOR2X1 U10208 ( .A(n16623), .B(n17114), .Y(n16778) );
  INVX1 U10209 ( .A(n17611), .Y(n16780) );
  NOR2X1 U10210 ( .A(n16780), .B(n17113), .Y(n16779) );
  BUFX2 U10211 ( .A(\lamb/scale_ls1/genblk1[1].mult/added[3] ), .Y(n16781) );
  BUFX2 U10212 ( .A(\lamb/scale_ls2/genblk1[0].mult/logB[2] ), .Y(n16782) );
  NOR2X1 U10213 ( .A(n16783), .B(n16784), .Y(n18365) );
  INVX1 U10214 ( .A(n18363), .Y(n16785) );
  INVX1 U10215 ( .A(n18364), .Y(n16786) );
  NOR2X1 U10216 ( .A(n16785), .B(n16786), .Y(n16783) );
  INVX1 U10217 ( .A(n18368), .Y(n16787) );
  INVX1 U10218 ( .A(n18370), .Y(n16788) );
  NOR2X1 U10219 ( .A(n16787), .B(n16788), .Y(n16784) );
  BUFX2 U10220 ( .A(n18602), .Y(n16789) );
  AND2X1 U10221 ( .A(n18674), .B(n18672), .Y(n18673) );
  INVX1 U10222 ( .A(n18673), .Y(n16790) );
  AND2X1 U10223 ( .A(n19302), .B(n19300), .Y(n19301) );
  INVX1 U10224 ( .A(n19301), .Y(n16791) );
  BUFX2 U10225 ( .A(n18662), .Y(n16792) );
  AND2X1 U10226 ( .A(n19340), .B(n19339), .Y(n19341) );
  INVX1 U10227 ( .A(n19341), .Y(n16793) );
  BUFX2 U10228 ( .A(n17892), .Y(n16794) );
  BUFX2 U10229 ( .A(n18451), .Y(n16795) );
  AND2X1 U10230 ( .A(n17985), .B(n17984), .Y(n17987) );
  INVX1 U10231 ( .A(n17987), .Y(n16796) );
  BUFX2 U10232 ( .A(n18743), .Y(n16797) );
  AND2X1 U10233 ( .A(n18612), .B(n18611), .Y(n18613) );
  INVX1 U10234 ( .A(n18613), .Y(n16798) );
  XOR2X1 U10235 ( .A(n18678), .B(n18694), .Y(n18612) );
  BUFX2 U10236 ( .A(n19126), .Y(n16799) );
  BUFX2 U10237 ( .A(n19056), .Y(n16800) );
  INVX1 U10238 ( .A(n16801), .Y(n17127) );
  INVX1 U10239 ( .A(n17330), .Y(n16802) );
  INVX1 U10240 ( .A(n17339), .Y(n16803) );
  NOR2X1 U10241 ( .A(n17336), .B(n16804), .Y(n16801) );
  NOR2X1 U10242 ( .A(n16802), .B(n16803), .Y(n16805) );
  INVX1 U10243 ( .A(n16805), .Y(n16804) );
  INVX1 U10244 ( .A(n18436), .Y(n16806) );
  AND2X1 U10245 ( .A(n19443), .B(n19486), .Y(n19446) );
  INVX1 U10246 ( .A(n19446), .Y(n16807) );
  AND2X1 U10247 ( .A(n16440), .B(n18472), .Y(n18473) );
  INVX1 U10248 ( .A(n18473), .Y(n16808) );
  INVX1 U10249 ( .A(n16809), .Y(n18463) );
  INVX1 U10250 ( .A(n18462), .Y(n16810) );
  INVX1 U10251 ( .A(n18535), .Y(n16811) );
  INVX1 U10252 ( .A(\lamb/scale_ls3/genblk1[1].mult/added[2] ), .Y(n16812) );
  NOR2X1 U10253 ( .A(n16812), .B(n16813), .Y(n16809) );
  NOR2X1 U10254 ( .A(n16810), .B(n16811), .Y(n16814) );
  INVX1 U10255 ( .A(n16814), .Y(n16813) );
  AND2X1 U10256 ( .A(n18152), .B(n16491), .Y(n18153) );
  INVX1 U10257 ( .A(n18153), .Y(n16815) );
  AND2X1 U10258 ( .A(n17980), .B(n16600), .Y(n17947) );
  INVX1 U10259 ( .A(n17947), .Y(n16816) );
  AND2X1 U10260 ( .A(\lamb/scale_ts1/genblk1[0].mult/added[2] ), .B(n17485), 
        .Y(n17472) );
  INVX1 U10261 ( .A(n17472), .Y(n16817) );
  BUFX2 U10262 ( .A(n18010), .Y(n16818) );
  AND2X1 U10263 ( .A(n18574), .B(n18485), .Y(n18480) );
  INVX1 U10264 ( .A(n18480), .Y(n16819) );
  AND2X1 U10265 ( .A(n18949), .B(n18811), .Y(n18814) );
  INVX1 U10266 ( .A(n18814), .Y(n16820) );
  BUFX2 U10267 ( .A(n17320), .Y(n16821) );
  AND2X1 U10268 ( .A(n17814), .B(n17819), .Y(n17818) );
  INVX1 U10269 ( .A(n17818), .Y(n16822) );
  INVX1 U10270 ( .A(n17847), .Y(n16823) );
  INVX1 U10271 ( .A(n16824), .Y(n18777) );
  INVX1 U10272 ( .A(n19259), .Y(n16825) );
  INVX1 U10273 ( .A(n18776), .Y(n16826) );
  INVX1 U10274 ( .A(n19569), .Y(n16827) );
  NOR2X1 U10275 ( .A(n16827), .B(n16828), .Y(n16824) );
  NOR2X1 U10276 ( .A(n16825), .B(n16826), .Y(n16829) );
  INVX1 U10277 ( .A(n16829), .Y(n16828) );
  AND2X1 U10278 ( .A(n16449), .B(n18775), .Y(n19569) );
  BUFX2 U10279 ( .A(n18043), .Y(n16830) );
  OR2X1 U10280 ( .A(n16774), .B(n16497), .Y(n17604) );
  INVX1 U10281 ( .A(n17604), .Y(n16831) );
  INVX1 U10282 ( .A(n16832), .Y(n18059) );
  INVX1 U10283 ( .A(n18057), .Y(n16833) );
  INVX1 U10284 ( .A(n18097), .Y(n16834) );
  INVX1 U10285 ( .A(n18058), .Y(n16835) );
  NOR2X1 U10286 ( .A(n16835), .B(n16836), .Y(n16832) );
  NOR2X1 U10287 ( .A(n16833), .B(n16834), .Y(n16837) );
  INVX1 U10288 ( .A(n16837), .Y(n16836) );
  BUFX2 U10289 ( .A(n17527), .Y(n16838) );
  OR2X1 U10290 ( .A(n17571), .B(n17574), .Y(n17524) );
  OR2X1 U10291 ( .A(n17614), .B(n17622), .Y(n17613) );
  INVX1 U10292 ( .A(n17613), .Y(n16839) );
  AND2X1 U10293 ( .A(n18458), .B(n18510), .Y(n18459) );
  INVX1 U10294 ( .A(n18459), .Y(n16840) );
  INVX1 U10295 ( .A(n16841), .Y(n17611) );
  INVX1 U10296 ( .A(n16392), .Y(n16842) );
  INVX1 U10297 ( .A(n18175), .Y(n16843) );
  NOR2X1 U10298 ( .A(n17610), .B(n16844), .Y(n16841) );
  NOR2X1 U10299 ( .A(n16842), .B(n16843), .Y(n16845) );
  INVX1 U10300 ( .A(n16845), .Y(n16844) );
  AND2X1 U10301 ( .A(n18587), .B(n18586), .Y(n18588) );
  BUFX2 U10302 ( .A(n18410), .Y(n16846) );
  NAND2X1 U10303 ( .A(n16847), .B(n16848), .Y(n18410) );
  INVX1 U10304 ( .A(n18408), .Y(n16849) );
  INVX1 U10305 ( .A(n18409), .Y(n16850) );
  NAND2X1 U10306 ( .A(n18531), .B(n16849), .Y(n16847) );
  NAND2X1 U10307 ( .A(n18531), .B(n16850), .Y(n16848) );
  INVX1 U10308 ( .A(n19174), .Y(n16851) );
  BUFX2 U10309 ( .A(\lamb/scale_ds3/genblk1[3].mult/logA[3] ), .Y(n16852) );
  NOR2X1 U10310 ( .A(n16853), .B(n16854), .Y(
        \lamb/scale_ds3/genblk1[3].mult/logA[3] ) );
  INVX1 U10311 ( .A(n17938), .Y(n16855) );
  INVX1 U10312 ( .A(n17939), .Y(n16856) );
  NOR2X1 U10313 ( .A(n16855), .B(n16856), .Y(n16853) );
  INVX1 U10314 ( .A(n17936), .Y(n16857) );
  INVX1 U10315 ( .A(n17937), .Y(n16858) );
  NOR2X1 U10316 ( .A(n16857), .B(n16858), .Y(n16854) );
  AND2X1 U10317 ( .A(n16622), .B(n16548), .Y(n17223) );
  INVX1 U10318 ( .A(n17223), .Y(n16859) );
  BUFX2 U10319 ( .A(\lamb/scale_ds2/genblk1[2].mult/logA[3] ), .Y(n16860) );
  NOR2X1 U10320 ( .A(n16861), .B(n16862), .Y(
        \lamb/scale_ds2/genblk1[2].mult/logA[3] ) );
  INVX1 U10321 ( .A(n18265), .Y(n16863) );
  INVX1 U10322 ( .A(n18266), .Y(n16864) );
  NOR2X1 U10323 ( .A(n16863), .B(n16864), .Y(n16861) );
  INVX1 U10324 ( .A(n18263), .Y(n16865) );
  INVX1 U10325 ( .A(n18264), .Y(n16866) );
  NOR2X1 U10326 ( .A(n16865), .B(n16866), .Y(n16862) );
  BUFX2 U10327 ( .A(n19584), .Y(n16867) );
  BUFX2 U10328 ( .A(n19550), .Y(n16868) );
  BUFX2 U10329 ( .A(n19109), .Y(n16869) );
  BUFX2 U10330 ( .A(n18505), .Y(n16870) );
  BUFX2 U10331 ( .A(n19108), .Y(n16871) );
  INVX1 U10332 ( .A(n16872), .Y(n19290) );
  INVX1 U10333 ( .A(n19287), .Y(n16873) );
  INVX1 U10334 ( .A(n19288), .Y(n16874) );
  NOR2X1 U10335 ( .A(n16618), .B(n16875), .Y(n16872) );
  NOR2X1 U10336 ( .A(n16873), .B(n16874), .Y(n16876) );
  INVX1 U10337 ( .A(n16876), .Y(n16875) );
  BUFX2 U10338 ( .A(n17878), .Y(n16877) );
  BUFX2 U10339 ( .A(n18143), .Y(n16878) );
  BUFX2 U10340 ( .A(n17787), .Y(n16879) );
  AND2X1 U10341 ( .A(n18369), .B(n17797), .Y(n17813) );
  INVX1 U10342 ( .A(n17813), .Y(n16880) );
  AND2X1 U10343 ( .A(n18099), .B(n18098), .Y(n18100) );
  INVX1 U10344 ( .A(n18100), .Y(n16881) );
  AND2X1 U10345 ( .A(\lamb/scale_ts0/genblk1[1].mult/added[2] ), .B(n17447), 
        .Y(n17423) );
  INVX1 U10346 ( .A(n17423), .Y(n16882) );
  AND2X1 U10347 ( .A(n19719), .B(n18349), .Y(n19720) );
  INVX1 U10348 ( .A(n19720), .Y(n16883) );
  AND2X1 U10349 ( .A(n18395), .B(n18394), .Y(n18542) );
  INVX1 U10350 ( .A(n18542), .Y(n16884) );
  AND2X1 U10351 ( .A(\lamb/scale_ls3/genblk1[2].mult/added[1] ), .B(n18477), 
        .Y(n18576) );
  INVX1 U10352 ( .A(n18576), .Y(n16885) );
  BUFX2 U10353 ( .A(n18352), .Y(n16886) );
  AND2X1 U10354 ( .A(n16566), .B(n18419), .Y(n18558) );
  INVX1 U10355 ( .A(n18558), .Y(n16887) );
  AND2X1 U10356 ( .A(n18029), .B(n18202), .Y(n18201) );
  INVX1 U10357 ( .A(n18201), .Y(n16888) );
  INVX1 U10358 ( .A(n19705), .Y(n16889) );
  AND2X1 U10359 ( .A(n16889), .B(n19704), .Y(n19707) );
  AND2X1 U10360 ( .A(n17941), .B(n17942), .Y(n17960) );
  INVX1 U10361 ( .A(n17960), .Y(n16890) );
  AND2X1 U10362 ( .A(n16890), .B(n17940), .Y(n17961) );
  AND2X1 U10363 ( .A(n17598), .B(n17601), .Y(n17581) );
  INVX1 U10364 ( .A(n17581), .Y(n16891) );
  AND2X1 U10365 ( .A(n19358), .B(n19357), .Y(n19369) );
  INVX1 U10366 ( .A(n19369), .Y(n16892) );
  AND2X1 U10367 ( .A(n16476), .B(n17125), .Y(n17323) );
  INVX1 U10368 ( .A(n17323), .Y(n16893) );
  AND2X1 U10369 ( .A(n16636), .B(n17541), .Y(n17559) );
  INVX1 U10370 ( .A(n17559), .Y(n16894) );
  OR2X1 U10371 ( .A(n17794), .B(n17793), .Y(n17831) );
  INVX1 U10372 ( .A(n17831), .Y(n16895) );
  AND2X1 U10373 ( .A(n18317), .B(n18316), .Y(n19739) );
  INVX1 U10374 ( .A(n19739), .Y(n16896) );
  AND2X1 U10375 ( .A(n18122), .B(n19772), .Y(n19700) );
  INVX1 U10376 ( .A(n19700), .Y(n16897) );
  AND2X1 U10377 ( .A(n18886), .B(n18866), .Y(n18856) );
  INVX1 U10378 ( .A(n18856), .Y(n16898) );
  AND2X1 U10379 ( .A(\lamb/scale_ds1/genblk1[3].mult/added[2] ), .B(n17316), 
        .Y(n17310) );
  INVX1 U10380 ( .A(n17310), .Y(n16899) );
  AND2X1 U10381 ( .A(n19272), .B(n18830), .Y(n18834) );
  INVX1 U10382 ( .A(n18834), .Y(n16900) );
  OR2X1 U10383 ( .A(n19267), .B(n16470), .Y(n18830) );
  AND2X1 U10384 ( .A(n18516), .B(n18402), .Y(n18465) );
  INVX1 U10385 ( .A(n18465), .Y(n16901) );
  OR2X1 U10386 ( .A(n19137), .B(n19136), .Y(n19170) );
  INVX1 U10387 ( .A(n19170), .Y(n16902) );
  AND2X1 U10388 ( .A(\lamb/scale_bs3/genblk1[1].mult/added[1] ), .B(n18470), 
        .Y(n18532) );
  INVX1 U10389 ( .A(n18532), .Y(n16903) );
  OR2X1 U10390 ( .A(n17589), .B(n17590), .Y(n17389) );
  INVX1 U10391 ( .A(n17389), .Y(n16904) );
  AND2X1 U10392 ( .A(n19418), .B(n19409), .Y(n19410) );
  INVX1 U10393 ( .A(n19410), .Y(n16905) );
  INVX1 U10394 ( .A(n17777), .Y(n16906) );
  INVX1 U10395 ( .A(n16907), .Y(n19319) );
  INVX1 U10396 ( .A(n19291), .Y(n16908) );
  INVX1 U10397 ( .A(n19292), .Y(n16909) );
  NOR2X1 U10398 ( .A(n19313), .B(n16910), .Y(n16907) );
  NOR2X1 U10399 ( .A(n16908), .B(n16909), .Y(n16911) );
  INVX1 U10400 ( .A(n16911), .Y(n16910) );
  BUFX2 U10401 ( .A(n18130), .Y(n16912) );
  BUFX2 U10402 ( .A(n19460), .Y(n16913) );
  AND2X1 U10403 ( .A(n18784), .B(n18927), .Y(n18807) );
  INVX1 U10404 ( .A(n18807), .Y(n16914) );
  INVX1 U10405 ( .A(n16915), .Y(n19322) );
  INVX1 U10406 ( .A(n19293), .Y(n16916) );
  INVX1 U10407 ( .A(n19294), .Y(n16917) );
  NOR2X1 U10408 ( .A(n19315), .B(n16918), .Y(n16915) );
  NOR2X1 U10409 ( .A(n16916), .B(n16917), .Y(n16919) );
  INVX1 U10410 ( .A(n16919), .Y(n16918) );
  AND2X1 U10411 ( .A(n16589), .B(n17857), .Y(n17875) );
  INVX1 U10412 ( .A(n17875), .Y(n16920) );
  AND2X1 U10413 ( .A(n18377), .B(n18378), .Y(n18750) );
  INVX1 U10414 ( .A(n18750), .Y(n16921) );
  BUFX2 U10415 ( .A(n17269), .Y(n16922) );
  OR2X1 U10416 ( .A(n19735), .B(n19734), .Y(n16312) );
  INVX1 U10417 ( .A(n16312), .Y(n16923) );
  BUFX2 U10418 ( .A(\lamb/scale_ts3/genblk1[2].mult/logA[2] ), .Y(n16924) );
  BUFX2 U10419 ( .A(\lamb/scale_ds2/genblk1[1].mult/logA[2] ), .Y(n16925) );
  AND2X1 U10420 ( .A(n18491), .B(n18431), .Y(n18553) );
  INVX1 U10421 ( .A(n18553), .Y(n16926) );
  BUFX2 U10422 ( .A(n18933), .Y(n16927) );
  AND2X1 U10423 ( .A(n18884), .B(n18874), .Y(n18868) );
  INVX1 U10424 ( .A(n18868), .Y(n16928) );
  AND2X1 U10425 ( .A(n19397), .B(n19415), .Y(n19436) );
  INVX1 U10426 ( .A(n19436), .Y(n16929) );
  INVX1 U10427 ( .A(n18897), .Y(n16930) );
  AND2X1 U10428 ( .A(n19079), .B(n19116), .Y(n19118) );
  INVX1 U10429 ( .A(n19118), .Y(n16931) );
  OR2X1 U10430 ( .A(n19081), .B(n19078), .Y(n19116) );
  INVX1 U10431 ( .A(n18294), .Y(n16932) );
  INVX1 U10432 ( .A(n16933), .Y(n17430) );
  INVX1 U10433 ( .A(n17394), .Y(n16934) );
  INVX1 U10434 ( .A(n17446), .Y(n16935) );
  NOR2X1 U10435 ( .A(n16935), .B(n16936), .Y(n16933) );
  NOR2X1 U10436 ( .A(n16934), .B(\lamb/scale_ts0/genblk1[1].mult/added[1] ), 
        .Y(n16937) );
  INVX1 U10437 ( .A(n16937), .Y(n16936) );
  BUFX2 U10438 ( .A(n19393), .Y(n16938) );
  AND2X1 U10439 ( .A(n18346), .B(n18345), .Y(n19718) );
  INVX1 U10440 ( .A(n19718), .Y(n16939) );
  AND2X1 U10441 ( .A(n18791), .B(n18934), .Y(n18901) );
  INVX1 U10442 ( .A(n18901), .Y(n16940) );
  AND2X1 U10443 ( .A(n18940), .B(n17073), .Y(n18934) );
  AND2X1 U10444 ( .A(\lamb/scale_ts1/genblk1[2].mult/added[1] ), .B(n17658), 
        .Y(n17697) );
  INVX1 U10445 ( .A(n17697), .Y(n16941) );
  BUFX2 U10446 ( .A(n17768), .Y(n16942) );
  NAND2X1 U10447 ( .A(n16943), .B(n16944), .Y(n17768) );
  INVX1 U10448 ( .A(n17763), .Y(n16945) );
  INVX1 U10449 ( .A(n16654), .Y(n16946) );
  INVX1 U10450 ( .A(n17764), .Y(n16947) );
  NAND2X1 U10451 ( .A(n16945), .B(n16946), .Y(n16943) );
  NAND2X1 U10452 ( .A(n16945), .B(n16947), .Y(n16944) );
  INVX1 U10453 ( .A(n16948), .Y(n18423) );
  INVX1 U10454 ( .A(n18416), .Y(n16949) );
  NOR2X1 U10455 ( .A(n16949), .B(n16950), .Y(n16948) );
  NOR2X1 U10456 ( .A(n18418), .B(\lamb/scale_bs3/genblk1[0].mult/added[1] ), 
        .Y(n16951) );
  INVX1 U10457 ( .A(n16951), .Y(n16950) );
  AND2X1 U10458 ( .A(n18786), .B(n16563), .Y(n18959) );
  INVX1 U10459 ( .A(n18959), .Y(n16952) );
  INVX1 U10460 ( .A(n16953), .Y(n19495) );
  INVX1 U10461 ( .A(n19472), .Y(n16954) );
  INVX1 U10462 ( .A(n19473), .Y(n16955) );
  INVX1 U10463 ( .A(n19493), .Y(n16956) );
  NOR2X1 U10464 ( .A(n16956), .B(n16957), .Y(n16953) );
  NOR2X1 U10465 ( .A(n16954), .B(n16955), .Y(n16958) );
  INVX1 U10466 ( .A(n16958), .Y(n16957) );
  AND2X1 U10467 ( .A(n16656), .B(n19157), .Y(n19183) );
  INVX1 U10468 ( .A(n19183), .Y(n16959) );
  OR2X1 U10469 ( .A(n17563), .B(n17561), .Y(n17565) );
  INVX1 U10470 ( .A(n17565), .Y(n16960) );
  OR2X1 U10471 ( .A(n17707), .B(\lamb/scale_ds1/genblk1[2].mult/added[2] ), 
        .Y(n17722) );
  INVX1 U10472 ( .A(n17722), .Y(n16961) );
  AND2X1 U10473 ( .A(\lamb/scale_bs2/genblk1[0].mult/added[3] ), .B(n17571), 
        .Y(n17530) );
  INVX1 U10474 ( .A(n17530), .Y(n16962) );
  AND2X1 U10475 ( .A(\lamb/scale_ts2/genblk1[3].mult/added[1] ), .B(n18071), 
        .Y(n18089) );
  INVX1 U10476 ( .A(n18089), .Y(n16963) );
  OR2X1 U10477 ( .A(\lamb/scale_ts3/genblk1[2].mult/added[1] ), .B(n18968), 
        .Y(n19006) );
  INVX1 U10478 ( .A(n19006), .Y(n16964) );
  AND2X1 U10479 ( .A(n19154), .B(n19156), .Y(n19160) );
  INVX1 U10480 ( .A(n19160), .Y(n16965) );
  AND2X1 U10481 ( .A(\lamb/scale_ts3/genblk1[3].mult/added[3] ), .B(n19127), 
        .Y(n19154) );
  BUFX2 U10482 ( .A(n17881), .Y(n16966) );
  BUFX2 U10483 ( .A(n17982), .Y(n16967) );
  INVX1 U10484 ( .A(n18270), .Y(n16968) );
  AND2X1 U10485 ( .A(n19360), .B(n19385), .Y(n19387) );
  INVX1 U10486 ( .A(n19387), .Y(n16969) );
  BUFX2 U10487 ( .A(n19013), .Y(n16970) );
  BUFX2 U10488 ( .A(n19492), .Y(n16971) );
  INVX1 U10489 ( .A(n16972), .Y(n17353) );
  INVX1 U10490 ( .A(n17328), .Y(n16973) );
  INVX1 U10491 ( .A(n17329), .Y(n16974) );
  INVX1 U10492 ( .A(\lamb/scale_ts1/genblk1[3].mult/added[1] ), .Y(n16975) );
  NOR2X1 U10493 ( .A(n16975), .B(n16976), .Y(n16972) );
  NOR2X1 U10494 ( .A(n16973), .B(n16974), .Y(n16977) );
  INVX1 U10495 ( .A(n16977), .Y(n16976) );
  AND2X1 U10496 ( .A(n17499), .B(n17502), .Y(n17497) );
  INVX1 U10497 ( .A(n17497), .Y(n16978) );
  AND2X1 U10498 ( .A(n16386), .B(n16978), .Y(n17500) );
  AND2X1 U10499 ( .A(n16623), .B(n18179), .Y(n19766) );
  INVX1 U10500 ( .A(n19766), .Y(n16979) );
  AND2X1 U10501 ( .A(n16404), .B(n16979), .Y(n19769) );
  AND2X1 U10502 ( .A(n19746), .B(n18314), .Y(n19738) );
  INVX1 U10503 ( .A(n19738), .Y(n16980) );
  INVX1 U10504 ( .A(n19266), .Y(n16981) );
  AND2X1 U10505 ( .A(n17596), .B(n17599), .Y(n18328) );
  INVX1 U10506 ( .A(n18328), .Y(n16982) );
  BUFX2 U10507 ( .A(n17375), .Y(n16983) );
  BUFX2 U10508 ( .A(n18075), .Y(n16984) );
  BUFX2 U10509 ( .A(n17734), .Y(n16985) );
  INVX1 U10510 ( .A(n18081), .Y(n16986) );
  AND2X1 U10511 ( .A(\lamb/scale_ds3/genblk1[2].mult/added[4] ), .B(
        \add_x_46/n1 ), .Y(n19020) );
  INVX1 U10512 ( .A(n19020), .Y(n16987) );
  AND2X1 U10513 ( .A(n16395), .B(n18430), .Y(n18548) );
  INVX1 U10514 ( .A(n18548), .Y(n16988) );
  BUFX2 U10515 ( .A(n17167), .Y(n16989) );
  BUFX2 U10516 ( .A(n17210), .Y(n16990) );
  BUFX2 U10517 ( .A(n19327), .Y(n16991) );
  NOR2X1 U10518 ( .A(n16992), .B(n16993), .Y(n19327) );
  INVX1 U10519 ( .A(n19271), .Y(n16994) );
  INVX1 U10520 ( .A(n19263), .Y(n16995) );
  NOR2X1 U10521 ( .A(n16994), .B(n16995), .Y(n16992) );
  INVX1 U10522 ( .A(n19261), .Y(n16996) );
  NOR2X1 U10523 ( .A(n16996), .B(n19262), .Y(n16993) );
  OR2X1 U10524 ( .A(n19260), .B(n19259), .Y(n19271) );
  AND2X1 U10525 ( .A(n17934), .B(n17925), .Y(n17926) );
  INVX1 U10526 ( .A(n17926), .Y(n16997) );
  INVX1 U10527 ( .A(n17836), .Y(n16998) );
  AND2X1 U10528 ( .A(n17670), .B(n17717), .Y(n17706) );
  INVX1 U10529 ( .A(n17706), .Y(n16999) );
  OR2X1 U10530 ( .A(n18260), .B(n18261), .Y(n18253) );
  INVX1 U10531 ( .A(n18253), .Y(n17000) );
  INVX1 U10532 ( .A(n18565), .Y(n17001) );
  AND2X1 U10533 ( .A(n18413), .B(n17666), .Y(n17340) );
  INVX1 U10534 ( .A(n17340), .Y(n17002) );
  AND2X1 U10535 ( .A(n16443), .B(n17623), .Y(n17644) );
  INVX1 U10536 ( .A(n17644), .Y(n17003) );
  AND2X1 U10537 ( .A(n18163), .B(n18160), .Y(n18170) );
  INVX1 U10538 ( .A(n18170), .Y(n17004) );
  AND2X1 U10539 ( .A(n19230), .B(n19225), .Y(n19221) );
  INVX1 U10540 ( .A(n19221), .Y(n17005) );
  AND2X1 U10541 ( .A(n18198), .B(n18206), .Y(n19661) );
  INVX1 U10542 ( .A(n19661), .Y(n17006) );
  AND2X1 U10543 ( .A(\add_x_52/n1 ), .B(
        \lamb/scale_ls3/genblk1[1].mult/added[4] ), .Y(n18455) );
  INVX1 U10544 ( .A(n18455), .Y(n17007) );
  AND2X1 U10545 ( .A(n19434), .B(n19433), .Y(n19432) );
  INVX1 U10546 ( .A(n19432), .Y(n17008) );
  INVX1 U10547 ( .A(n17989), .Y(n17009) );
  BUFX2 U10548 ( .A(n17806), .Y(n17010) );
  AND2X1 U10549 ( .A(n16527), .B(n19250), .Y(n19514) );
  INVX1 U10550 ( .A(n19514), .Y(n17011) );
  AND2X1 U10551 ( .A(\lamb/scale_ls2/genblk1[2].mult/added[4] ), .B(
        \add_x_64/n1 ), .Y(n18114) );
  INVX1 U10552 ( .A(n18114), .Y(n17012) );
  AND2X1 U10553 ( .A(\lamb/scale_ls2/genblk1[1].mult/added[3] ), .B(n18117), 
        .Y(n18128) );
  INVX1 U10554 ( .A(n18128), .Y(n17013) );
  AND2X1 U10555 ( .A(n18974), .B(n18975), .Y(n19023) );
  INVX1 U10556 ( .A(n19023), .Y(n17014) );
  AND2X1 U10557 ( .A(n17654), .B(n16509), .Y(n17701) );
  INVX1 U10558 ( .A(n17701), .Y(n17015) );
  AND2X1 U10559 ( .A(n17481), .B(n17480), .Y(n18267) );
  INVX1 U10560 ( .A(n18267), .Y(n17016) );
  AND2X1 U10561 ( .A(n18268), .B(n17016), .Y(n18274) );
  AND2X1 U10562 ( .A(\lamb/scale_ts1/genblk1[1].mult/added[2] ), .B(n16945), 
        .Y(n17820) );
  INVX1 U10563 ( .A(n17820), .Y(n17017) );
  INVX1 U10564 ( .A(n17755), .Y(n17018) );
  AND2X1 U10565 ( .A(n16524), .B(n17407), .Y(n17449) );
  INVX1 U10566 ( .A(n17449), .Y(n17019) );
  BUFX2 U10567 ( .A(n18371), .Y(n17020) );
  AND2X1 U10568 ( .A(n16810), .B(n16812), .Y(n18534) );
  INVX1 U10569 ( .A(n18534), .Y(n17021) );
  AND2X1 U10570 ( .A(n18336), .B(n18335), .Y(n19664) );
  INVX1 U10571 ( .A(n19664), .Y(n17022) );
  INVX1 U10572 ( .A(n19334), .Y(n17023) );
  OR2X1 U10573 ( .A(n18234), .B(n18233), .Y(n18232) );
  INVX1 U10574 ( .A(n18232), .Y(n17024) );
  BUFX2 U10575 ( .A(n17275), .Y(n17025) );
  OR2X1 U10576 ( .A(n18382), .B(n18380), .Y(n18388) );
  INVX1 U10577 ( .A(n18388), .Y(n17026) );
  INVX1 U10578 ( .A(n19146), .Y(n17027) );
  BUFX2 U10579 ( .A(\lamb/scale_ts0/genblk1[0].mult/logA[1] ), .Y(n17028) );
  AND2X1 U10580 ( .A(n18242), .B(n18241), .Y(n19757) );
  INVX1 U10581 ( .A(n19757), .Y(n17029) );
  BUFX2 U10582 ( .A(n17233), .Y(n17030) );
  OR2X1 U10583 ( .A(n18301), .B(n18752), .Y(n16307) );
  INVX1 U10584 ( .A(n16307), .Y(n17031) );
  AND2X1 U10585 ( .A(n19750), .B(n19749), .Y(n17723) );
  INVX1 U10586 ( .A(n17723), .Y(n17032) );
  AND2X1 U10587 ( .A(n18985), .B(n18984), .Y(n19025) );
  INVX1 U10588 ( .A(n19025), .Y(n17033) );
  AND2X1 U10589 ( .A(\lamb/scale_bs3/genblk1[1].mult/added[3] ), .B(n18397), 
        .Y(n18526) );
  INVX1 U10590 ( .A(n18526), .Y(n17034) );
  INVX1 U10591 ( .A(n17362), .Y(n17035) );
  AND2X1 U10592 ( .A(n19699), .B(n18342), .Y(n19666) );
  AND2X1 U10593 ( .A(n17515), .B(n17513), .Y(n17522) );
  INVX1 U10594 ( .A(n17522), .Y(n17036) );
  BUFX2 U10595 ( .A(n19683), .Y(n17037) );
  BUFX2 U10596 ( .A(n17221), .Y(n17038) );
  BUFX2 U10597 ( .A(n17374), .Y(n17039) );
  AND2X1 U10598 ( .A(n17627), .B(n17626), .Y(n18356) );
  INVX1 U10599 ( .A(n18356), .Y(n17040) );
  OR2X1 U10600 ( .A(\lamb/scale_ds2/genblk1[3].mult/added[4] ), .B(
        \add_x_58/n1 ), .Y(n18038) );
  INVX1 U10601 ( .A(n18038), .Y(n17041) );
  AND2X1 U10602 ( .A(\lamb/scale_ds1/genblk1[1].mult/added[4] ), .B(
        \add_x_73/n1 ), .Y(n17776) );
  INVX1 U10603 ( .A(n17776), .Y(n17042) );
  BUFX2 U10604 ( .A(n19275), .Y(n17043) );
  AND2X1 U10605 ( .A(\lamb/scale_ls3/genblk1[0].mult/added[2] ), .B(
        \lamb/scale_ls3/genblk1[0].mult/added[1] ), .Y(n18550) );
  INVX1 U10606 ( .A(n18550), .Y(n17044) );
  AND2X1 U10607 ( .A(\lamb/scale_ds2/genblk1[1].mult/added[4] ), .B(
        \add_x_60/n1 ), .Y(n17965) );
  INVX1 U10608 ( .A(n17965), .Y(n17045) );
  BUFX2 U10609 ( .A(n18848), .Y(n17046) );
  AND2X1 U10610 ( .A(n18337), .B(n18334), .Y(n19697) );
  INVX1 U10611 ( .A(n19697), .Y(n17047) );
  AND2X1 U10612 ( .A(\lamb/scale_ts2/genblk1[3].mult/added[3] ), .B(n18025), 
        .Y(n18078) );
  INVX1 U10613 ( .A(n18078), .Y(n17048) );
  BUFX2 U10614 ( .A(n19675), .Y(n17049) );
  AND2X1 U10615 ( .A(\lamb/scale_ts2/genblk1[2].mult/added[3] ), .B(n17870), 
        .Y(n17911) );
  INVX1 U10616 ( .A(n17911), .Y(n17050) );
  AND2X1 U10617 ( .A(n19594), .B(n16736), .Y(n19519) );
  INVX1 U10618 ( .A(n19519), .Y(n17051) );
  BUFX2 U10619 ( .A(n17533), .Y(n17052) );
  BUFX2 U10620 ( .A(n19033), .Y(n17053) );
  AND2X1 U10621 ( .A(n16446), .B(n18507), .Y(n18513) );
  INVX1 U10622 ( .A(n18513), .Y(n17054) );
  AND2X1 U10623 ( .A(n17054), .B(n18461), .Y(n18535) );
  AND2X1 U10624 ( .A(n19052), .B(n19039), .Y(n19069) );
  INVX1 U10625 ( .A(n19069), .Y(n17055) );
  BUFX2 U10626 ( .A(n19311), .Y(n17056) );
  NOR2X1 U10627 ( .A(n17057), .B(n17058), .Y(n19311) );
  INVX1 U10628 ( .A(n19270), .Y(n17059) );
  NOR2X1 U10629 ( .A(n19271), .B(n17059), .Y(n17057) );
  INVX1 U10630 ( .A(n19268), .Y(n17060) );
  NOR2X1 U10631 ( .A(n17060), .B(n19269), .Y(n17058) );
  AND2X1 U10632 ( .A(n16723), .B(n16413), .Y(n19268) );
  BUFX2 U10633 ( .A(n19475), .Y(n17061) );
  AND2X1 U10634 ( .A(n18245), .B(n19762), .Y(n19761) );
  INVX1 U10635 ( .A(n19761), .Y(n17062) );
  AND2X1 U10636 ( .A(n16530), .B(n17864), .Y(n17903) );
  INVX1 U10637 ( .A(n17903), .Y(n17063) );
  BUFX2 U10638 ( .A(n19346), .Y(n17064) );
  AND2X1 U10639 ( .A(\lamb/scale_ds1/genblk1[3].mult/added[4] ), .B(
        \add_x_71/n1 ), .Y(n17343) );
  INVX1 U10640 ( .A(n17343), .Y(n17065) );
  INVX1 U10641 ( .A(n18833), .Y(n17066) );
  OR2X1 U10642 ( .A(n17256), .B(n17255), .Y(n17299) );
  INVX1 U10643 ( .A(n17299), .Y(n17067) );
  BUFX2 U10644 ( .A(\lamb/scale_ts0/genblk1[2].mult/logA[1] ), .Y(n17068) );
  OR2X1 U10645 ( .A(n16580), .B(n19622), .Y(n19578) );
  INVX1 U10646 ( .A(n19578), .Y(n17069) );
  OR2X1 U10647 ( .A(n19082), .B(n19356), .Y(n19178) );
  INVX1 U10648 ( .A(n19178), .Y(n17070) );
  AND2X1 U10649 ( .A(n16494), .B(n19241), .Y(n19456) );
  INVX1 U10650 ( .A(n19456), .Y(n17071) );
  AND2X1 U10651 ( .A(n16551), .B(n18825), .Y(n18655) );
  INVX1 U10652 ( .A(n18655), .Y(n17072) );
  BUFX2 U10653 ( .A(n18941), .Y(n17073) );
  AND2X1 U10654 ( .A(n18906), .B(n18768), .Y(n18923) );
  INVX1 U10655 ( .A(n18923), .Y(n17074) );
  BUFX2 U10656 ( .A(n18288), .Y(n17075) );
  BUFX2 U10657 ( .A(n19238), .Y(n17076) );
  BUFX2 U10658 ( .A(n19065), .Y(n17077) );
  INVX1 U10659 ( .A(n18769), .Y(n17078) );
  OR2X1 U10660 ( .A(n18747), .B(n17078), .Y(n18816) );
  BUFX2 U10661 ( .A(n19756), .Y(n17079) );
  BUFX2 U10662 ( .A(n19708), .Y(n17080) );
  BUFX2 U10663 ( .A(n17460), .Y(n17081) );
  BUFX2 U10664 ( .A(n17181), .Y(n17082) );
  AND2X1 U10665 ( .A(\add_x_45/n1 ), .B(n19100), .Y(n19164) );
  INVX1 U10666 ( .A(n19164), .Y(n17083) );
  BUFX2 U10667 ( .A(\lamb/scale_bs3/genblk1[0].mult/logB[3] ), .Y(n17084) );
  BUFX2 U10668 ( .A(\lamb/scale_bs2/genblk1[1].mult/added[4] ), .Y(n17085) );
  NOR2X1 U10669 ( .A(n17086), .B(n17087), .Y(
        \lamb/scale_bs2/genblk1[1].mult/added[4] ) );
  INVX1 U10670 ( .A(n19716), .Y(n17088) );
  INVX1 U10671 ( .A(n19773), .Y(n17089) );
  NOR2X1 U10672 ( .A(n17088), .B(n17089), .Y(n17086) );
  INVX1 U10673 ( .A(n19714), .Y(n17090) );
  INVX1 U10674 ( .A(n19715), .Y(n17091) );
  NOR2X1 U10675 ( .A(n17090), .B(n17091), .Y(n17087) );
  INVX1 U10676 ( .A(n18875), .Y(n17092) );
  BUFX2 U10677 ( .A(n17270), .Y(n17093) );
  BUFX2 U10678 ( .A(n17751), .Y(n17094) );
  OR2X1 U10679 ( .A(\lamb/scale_ts0/genblk1[2].mult/added[4] ), .B(
        \add_x_77/n1 ), .Y(n17264) );
  INVX1 U10680 ( .A(n17264), .Y(n17095) );
  BUFX2 U10681 ( .A(n19592), .Y(n17096) );
  NAND2X1 U10682 ( .A(n17097), .B(n17098), .Y(n19592) );
  INVX1 U10683 ( .A(n18756), .Y(n17099) );
  INVX1 U10684 ( .A(n16506), .Y(n17100) );
  INVX1 U10685 ( .A(n18760), .Y(n17101) );
  NAND2X1 U10686 ( .A(n17099), .B(n17100), .Y(n17097) );
  NAND2X1 U10687 ( .A(n17099), .B(n17101), .Y(n17098) );
  BUFX2 U10688 ( .A(n18197), .Y(n17102) );
  INVX1 U10689 ( .A(n19544), .Y(n17103) );
  BUFX2 U10690 ( .A(\lamb/scale_bs3/genblk1[0].mult/logB[1] ), .Y(n17104) );
  BUFX2 U10691 ( .A(\lamb/scale_bs2/genblk1[1].mult/added[2] ), .Y(n17105) );
  BUFX2 U10692 ( .A(\lamb/scale_ts1/genblk1[0].mult/logB[2] ), .Y(n17106) );
  AND2X1 U10693 ( .A(n16762), .B(n18908), .Y(n18952) );
  INVX1 U10694 ( .A(n18952), .Y(n17107) );
  AND2X1 U10695 ( .A(n18490), .B(n18573), .Y(n18717) );
  INVX1 U10696 ( .A(n18717), .Y(n17108) );
  BUFX2 U10697 ( .A(\lamb/scale_ls3/genblk1[0].mult/logB[2] ), .Y(n17109) );
  NAND2X1 U10698 ( .A(n17110), .B(n17111), .Y(
        \lamb/scale_ls3/genblk1[0].mult/logB[2] ) );
  INVX1 U10699 ( .A(n18177), .Y(n17112) );
  INVX1 U10700 ( .A(n18178), .Y(n17113) );
  INVX1 U10701 ( .A(n16617), .Y(n17114) );
  NAND2X1 U10702 ( .A(n17112), .B(n17113), .Y(n17110) );
  NAND2X1 U10703 ( .A(n17112), .B(n17114), .Y(n17111) );
  INVX1 U10704 ( .A(n18720), .Y(n17115) );
  AND2X1 U10705 ( .A(n16533), .B(n18573), .Y(n18685) );
  INVX1 U10706 ( .A(n18685), .Y(n17116) );
  BUFX2 U10707 ( .A(n16313), .Y(n17117) );
  NOR2X1 U10708 ( .A(n17118), .B(n17119), .Y(n16313) );
  INVX1 U10709 ( .A(n19730), .Y(n17120) );
  NOR2X1 U10710 ( .A(n17120), .B(n16733), .Y(n17118) );
  INVX1 U10711 ( .A(n19728), .Y(n17121) );
  INVX1 U10712 ( .A(n19729), .Y(n17122) );
  NOR2X1 U10713 ( .A(n17121), .B(n17122), .Y(n17119) );
  AND2X1 U10714 ( .A(n17597), .B(n17605), .Y(n18156) );
  INVX1 U10715 ( .A(n18156), .Y(n17123) );
  BUFX2 U10716 ( .A(\lamb/scale_ls1/genblk1[1].mult/added[2] ), .Y(n17124) );
  OR2X1 U10717 ( .A(\lamb/scale_ts1/genblk1[3].mult/added[4] ), .B(
        \add_x_67/n1 ), .Y(n17324) );
  AOI21X1 U10718 ( .A(\add_x_67/n1 ), .B(
        \lamb/scale_ts1/genblk1[3].mult/added[4] ), .C(
        \lamb/scale_ts1/genblk1[3].mult/added[3] ), .Y(n17325) );
  INVX1 U10719 ( .A(n17325), .Y(n17125) );
  NOR3X1 U10720 ( .A(\lamb/scale_ts1/genblk1[3].mult/added[4] ), .B(
        \add_x_67/n1 ), .C(\lamb/scale_ts1/genblk1[3].mult/added[3] ), .Y(
        n17336) );
  NAND3X1 U10721 ( .A(\lamb/scale_ts1/genblk1[3].mult/added[4] ), .B(
        \add_x_67/n1 ), .C(\lamb/scale_ts1/genblk1[3].mult/added[3] ), .Y(
        n17128) );
  NAND3X1 U10722 ( .A(\lamb/scale_ts1/genblk1[3].mult/added[2] ), .B(
        \lamb/scale_ts1/genblk1[3].mult/added[1] ), .C(n17128), .Y(n17339) );
  NOR2X1 U10723 ( .A(\lamb/scale_ts1/genblk1[3].mult/added[1] ), .B(n16476), 
        .Y(n17130) );
  NAND2X1 U10724 ( .A(\lamb/scale_ts1/genblk1[3].mult/added[4] ), .B(
        \add_x_67/n1 ), .Y(n17129) );
  INVX1 U10725 ( .A(n17129), .Y(n17126) );
  NAND2X1 U10726 ( .A(\lamb/scale_ts1/genblk1[3].mult/added[2] ), .B(n17338), 
        .Y(n17329) );
  NAND3X1 U10727 ( .A(n17130), .B(n17126), .C(n16974), .Y(n17330) );
  AOI21X1 U10728 ( .A(\lamb/scale_ts1/genblk1[3].mult/added[1] ), .B(n17323), 
        .C(n17127), .Y(n17224) );
  INVX1 U10729 ( .A(n17128), .Y(n17132) );
  NAND2X1 U10730 ( .A(n17130), .B(n17129), .Y(n17355) );
  NAND3X1 U10731 ( .A(\lamb/scale_ts1/genblk1[3].mult/added[2] ), .B(n17355), 
        .C(n17338), .Y(n17131) );
  OAI21X1 U10732 ( .A(\lamb/scale_ts1/genblk1[3].mult/added[2] ), .B(n17132), 
        .C(n17131), .Y(n17342) );
  INVX1 U10733 ( .A(msg[47]), .Y(n17166) );
  INVX1 U10734 ( .A(msg[31]), .Y(n19551) );
  INVX1 U10735 ( .A(msg[3]), .Y(n19643) );
  AOI22X1 U10736 ( .A(msg[3]), .B(msg[31]), .C(n19551), .D(n19643), .Y(n19683)
         );
  MUX2X1 U10737 ( .B(n17166), .A(msg[47]), .S(n17037), .Y(n17433) );
  INVX1 U10738 ( .A(msg[39]), .Y(n19525) );
  INVX1 U10739 ( .A(msg[51]), .Y(n17457) );
  INVX1 U10740 ( .A(msg[15]), .Y(n19597) );
  INVX1 U10741 ( .A(msg[35]), .Y(n19536) );
  MUX2X1 U10742 ( .B(msg[15]), .A(n19597), .S(n19536), .Y(n17215) );
  MUX2X1 U10743 ( .B(n17457), .A(msg[51]), .S(n17215), .Y(n17432) );
  MUX2X1 U10744 ( .B(n19525), .A(msg[39]), .S(n17432), .Y(n17293) );
  INVX1 U10745 ( .A(msg[23]), .Y(n19572) );
  INVX1 U10746 ( .A(msg[43]), .Y(n19450) );
  AOI22X1 U10747 ( .A(msg[43]), .B(msg[23]), .C(n19572), .D(n19450), .Y(n17135) );
  INVX1 U10748 ( .A(msg[59]), .Y(n19668) );
  INVX1 U10749 ( .A(msg[11]), .Y(n19609) );
  INVX1 U10750 ( .A(msg[19]), .Y(n19583) );
  INVX1 U10751 ( .A(msg[7]), .Y(n19626) );
  INVX1 U10752 ( .A(msg[27]), .Y(n19561) );
  MUX2X1 U10753 ( .B(msg[7]), .A(n19626), .S(n19561), .Y(n19682) );
  MUX2X1 U10754 ( .B(n19583), .A(msg[19]), .S(n19682), .Y(n17162) );
  MUX2X1 U10755 ( .B(n19609), .A(msg[11]), .S(n17162), .Y(n17133) );
  MUX2X1 U10756 ( .B(msg[59]), .A(n19668), .S(n17133), .Y(n17134) );
  FAX1 U10757 ( .A(msg[55]), .B(n16667), .C(n17134), .YS(n17136) );
  FAX1 U10758 ( .A(n17433), .B(n17293), .C(n17136), .YS(n17222) );
  INVX1 U10759 ( .A(msg[45]), .Y(n17376) );
  INVX1 U10760 ( .A(msg[21]), .Y(n19576) );
  INVX1 U10761 ( .A(msg[41]), .Y(n19509) );
  AOI22X1 U10762 ( .A(msg[41]), .B(msg[21]), .C(n19576), .D(n19509), .Y(n17167) );
  MUX2X1 U10763 ( .B(n17376), .A(msg[45]), .S(n16989), .Y(n17155) );
  INVX1 U10764 ( .A(msg[25]), .Y(n19565) );
  INVX1 U10765 ( .A(msg[33]), .Y(n19669) );
  INVX1 U10766 ( .A(msg[13]), .Y(n19601) );
  INVX1 U10767 ( .A(msg[1]), .Y(n19651) );
  AOI22X1 U10768 ( .A(msg[1]), .B(msg[13]), .C(n19601), .D(n19651), .Y(n17137)
         );
  MUX2X1 U10769 ( .B(n19669), .A(msg[33]), .S(n17137), .Y(n17138) );
  MUX2X1 U10770 ( .B(n19565), .A(msg[25]), .S(n17138), .Y(n17143) );
  INVX1 U10771 ( .A(msg[9]), .Y(n19615) );
  INVX1 U10772 ( .A(msg[29]), .Y(n19555) );
  MUX2X1 U10773 ( .B(msg[9]), .A(n19615), .S(n19555), .Y(n17246) );
  INVX1 U10774 ( .A(msg[17]), .Y(n19587) );
  INVX1 U10775 ( .A(msg[37]), .Y(n19529) );
  MUX2X1 U10776 ( .B(msg[17]), .A(n19587), .S(n19529), .Y(n17254) );
  INVX1 U10777 ( .A(msg[57]), .Y(n17199) );
  INVX1 U10778 ( .A(msg[5]), .Y(n19632) );
  INVX1 U10779 ( .A(msg[53]), .Y(n17283) );
  INVX1 U10780 ( .A(msg[49]), .Y(n17187) );
  MUX2X1 U10781 ( .B(msg[53]), .A(n17283), .S(n17187), .Y(n17139) );
  MUX2X1 U10782 ( .B(n19632), .A(msg[5]), .S(n17139), .Y(n17140) );
  MUX2X1 U10783 ( .B(msg[57]), .A(n17199), .S(n17140), .Y(n17141) );
  FAX1 U10784 ( .A(n17246), .B(n17254), .C(n17141), .YS(n17142) );
  FAX1 U10785 ( .A(n17155), .B(n17143), .C(n17142), .YS(n17588) );
  INVX1 U10786 ( .A(msg[18]), .Y(n19585) );
  INVX1 U10787 ( .A(msg[38]), .Y(n19527) );
  MUX2X1 U10788 ( .B(msg[18]), .A(n19585), .S(n19527), .Y(n17165) );
  INVX1 U10789 ( .A(msg[30]), .Y(n19553) );
  MUX2X1 U10790 ( .B(n19553), .A(msg[30]), .S(msg[54]), .Y(n17399) );
  INVX1 U10791 ( .A(msg[46]), .Y(n17185) );
  INVX1 U10792 ( .A(msg[42]), .Y(n19670) );
  INVX1 U10793 ( .A(msg[22]), .Y(n19574) );
  AOI22X1 U10794 ( .A(msg[22]), .B(msg[42]), .C(n19670), .D(n19574), .Y(n17181) );
  MUX2X1 U10795 ( .B(n17185), .A(msg[46]), .S(n17082), .Y(n17248) );
  INVX1 U10796 ( .A(msg[2]), .Y(n19647) );
  INVX1 U10797 ( .A(msg[26]), .Y(n19563) );
  INVX1 U10798 ( .A(msg[6]), .Y(n19629) );
  AOI22X1 U10799 ( .A(msg[6]), .B(msg[26]), .C(n19563), .D(n19629), .Y(n17144)
         );
  MUX2X1 U10800 ( .B(n19647), .A(msg[2]), .S(n17144), .Y(n17145) );
  FAX1 U10801 ( .A(n17248), .B(msg[58]), .C(n17145), .YS(n17146) );
  FAX1 U10802 ( .A(n17165), .B(n17399), .C(n17146), .YS(n17148) );
  INVX1 U10803 ( .A(msg[14]), .Y(n19599) );
  INVX1 U10804 ( .A(msg[34]), .Y(n19539) );
  MUX2X1 U10805 ( .B(msg[14]), .A(n19599), .S(n19539), .Y(n17285) );
  INVX1 U10806 ( .A(n17285), .Y(n17211) );
  INVX1 U10807 ( .A(msg[10]), .Y(n19612) );
  MUX2X1 U10808 ( .B(n19612), .A(msg[10]), .S(msg[50]), .Y(n17412) );
  INVX1 U10809 ( .A(n17412), .Y(n17147) );
  FAX1 U10810 ( .A(n17148), .B(n17211), .C(n17147), .YS(n17578) );
  INVX1 U10811 ( .A(msg[32]), .Y(n19546) );
  INVX1 U10812 ( .A(msg[24]), .Y(n19568) );
  INVX1 U10813 ( .A(msg[4]), .Y(n19637) );
  AOI22X1 U10814 ( .A(msg[4]), .B(n19568), .C(msg[24]), .D(n19637), .Y(n17398)
         );
  MUX2X1 U10815 ( .B(msg[32]), .A(n19546), .S(n16591), .Y(n17288) );
  INVX1 U10816 ( .A(msg[0]), .Y(n19656) );
  INVX1 U10817 ( .A(msg[16]), .Y(n19590) );
  INVX1 U10818 ( .A(msg[36]), .Y(n19533) );
  MUX2X1 U10819 ( .B(msg[16]), .A(n19590), .S(n19533), .Y(n17274) );
  MUX2X1 U10820 ( .B(n19656), .A(msg[0]), .S(n17274), .Y(n17153) );
  INVX1 U10821 ( .A(msg[48]), .Y(n17290) );
  INVX1 U10822 ( .A(msg[44]), .Y(n19671) );
  MUX2X1 U10823 ( .B(msg[48]), .A(n17290), .S(n19671), .Y(n17411) );
  INVX1 U10824 ( .A(msg[40]), .Y(n19522) );
  INVX1 U10825 ( .A(msg[8]), .Y(n19619) );
  AOI22X1 U10826 ( .A(msg[8]), .B(msg[40]), .C(n19522), .D(n19619), .Y(n17151)
         );
  INVX1 U10827 ( .A(msg[20]), .Y(n19580) );
  INVX1 U10828 ( .A(msg[56]), .Y(n17231) );
  INVX1 U10829 ( .A(msg[28]), .Y(n19559) );
  INVX1 U10830 ( .A(msg[12]), .Y(n19605) );
  INVX1 U10831 ( .A(msg[52]), .Y(n17213) );
  AOI22X1 U10832 ( .A(msg[52]), .B(msg[12]), .C(n19605), .D(n17213), .Y(n17460) );
  MUX2X1 U10833 ( .B(n19559), .A(msg[28]), .S(n17081), .Y(n17439) );
  MUX2X1 U10834 ( .B(n17231), .A(msg[56]), .S(n17439), .Y(n17149) );
  MUX2X1 U10835 ( .B(msg[20]), .A(n19580), .S(n17149), .Y(n17150) );
  FAX1 U10836 ( .A(n17411), .B(n16668), .C(n17150), .YS(n17152) );
  FAX1 U10837 ( .A(n17288), .B(n17153), .C(n17152), .YS(n17579) );
  NAND2X1 U10838 ( .A(n16642), .B(n17579), .Y(n17154) );
  OR2X1 U10839 ( .A(n16548), .B(n17154), .Y(n17630) );
  AOI22X1 U10840 ( .A(msg[11]), .B(msg[13]), .C(n19601), .D(n19609), .Y(n19675) );
  MUX2X1 U10841 ( .B(n19565), .A(msg[25]), .S(n17049), .Y(n17175) );
  FAX1 U10842 ( .A(n17155), .B(msg[17]), .C(n17175), .YS(n17209) );
  MUX2X1 U10843 ( .B(n19553), .A(msg[30]), .S(n17274), .Y(n17291) );
  FAX1 U10844 ( .A(n17082), .B(n17165), .C(n17291), .YS(n17164) );
  AOI22X1 U10845 ( .A(msg[14]), .B(msg[28]), .C(n19559), .D(n19599), .Y(n17158) );
  AOI22X1 U10846 ( .A(msg[57]), .B(msg[10]), .C(n19612), .D(n17199), .Y(n17157) );
  AOI22X1 U10847 ( .A(msg[39]), .B(msg[33]), .C(n19669), .D(n19525), .Y(n17374) );
  MUX2X1 U10848 ( .B(n19580), .A(msg[20]), .S(msg[54]), .Y(n17234) );
  HAX1 U10849 ( .A(n17039), .B(n17234), .YS(n17156) );
  FAX1 U10850 ( .A(n16711), .B(n16669), .C(n17156), .YS(n17161) );
  HAX1 U10851 ( .A(n17432), .B(n17411), .YS(n17251) );
  MUX2X1 U10852 ( .B(n19656), .A(msg[0]), .S(n17251), .Y(n17159) );
  MUX2X1 U10853 ( .B(msg[24]), .A(n19568), .S(n17159), .Y(n17160) );
  FAX1 U10854 ( .A(n17162), .B(n17161), .C(n17160), .YS(n17163) );
  FAX1 U10855 ( .A(n17209), .B(n17164), .C(n17163), .YS(n17739) );
  INVX1 U10856 ( .A(n17739), .Y(n17589) );
  MUX2X1 U10857 ( .B(n19551), .A(msg[31]), .S(n17254), .Y(n17183) );
  MUX2X1 U10858 ( .B(n17166), .A(msg[47]), .S(n17165), .Y(n17418) );
  AOI22X1 U10859 ( .A(msg[3]), .B(msg[6]), .C(n19629), .D(n19643), .Y(n17284)
         );
  MUX2X1 U10860 ( .B(msg[9]), .A(n19615), .S(n16714), .Y(n17381) );
  INVX1 U10861 ( .A(n17381), .Y(n17382) );
  HAX1 U10862 ( .A(n16989), .B(n17412), .YS(n17435) );
  HAX1 U10863 ( .A(n17382), .B(n17435), .YS(n17217) );
  MUX2X1 U10864 ( .B(n17283), .A(msg[53]), .S(n17049), .Y(n17220) );
  MUX2X1 U10865 ( .B(n19568), .A(msg[24]), .S(n17220), .Y(n17250) );
  MUX2X1 U10866 ( .B(msg[20]), .A(n19580), .S(n17211), .Y(n17194) );
  MUX2X1 U10867 ( .B(n19522), .A(msg[40]), .S(n17215), .Y(n17236) );
  MUX2X1 U10868 ( .B(n17231), .A(msg[56]), .S(n17236), .Y(n17168) );
  MUX2X1 U10869 ( .B(n19590), .A(msg[16]), .S(n17168), .Y(n17169) );
  MUX2X1 U10870 ( .B(n19626), .A(msg[7]), .S(n17169), .Y(n17172) );
  AOI22X1 U10871 ( .A(msg[23]), .B(msg[26]), .C(n19563), .D(n19572), .Y(n17191) );
  MUX2X1 U10872 ( .B(msg[29]), .A(n19555), .S(n16592), .Y(n17379) );
  MUX2X1 U10873 ( .B(msg[44]), .A(n19671), .S(n17379), .Y(n17462) );
  MUX2X1 U10874 ( .B(n19605), .A(msg[12]), .S(n17462), .Y(n17170) );
  MUX2X1 U10875 ( .B(msg[32]), .A(n19546), .S(n17170), .Y(n17171) );
  FAX1 U10876 ( .A(n17194), .B(n17172), .C(n17171), .YS(n17173) );
  FAX1 U10877 ( .A(n17217), .B(n17250), .C(n17173), .YS(n17174) );
  FAX1 U10878 ( .A(n17183), .B(n17418), .C(n17174), .YS(n17716) );
  INVX1 U10879 ( .A(n17716), .Y(n17590) );
  HAX1 U10880 ( .A(n17439), .B(n17194), .YS(n17280) );
  MUX2X1 U10881 ( .B(msg[33]), .A(n19669), .S(n17185), .Y(n17192) );
  MUX2X1 U10882 ( .B(n19647), .A(msg[2]), .S(n17192), .Y(n17200) );
  HAX1 U10883 ( .A(n17200), .B(n17183), .YS(n17292) );
  MUX2X1 U10884 ( .B(msg[49]), .A(n17187), .S(n17381), .Y(n17273) );
  FAX1 U10885 ( .A(n17292), .B(n17273), .C(n17175), .YS(n17463) );
  AOI22X1 U10886 ( .A(msg[59]), .B(msg[10]), .C(n19612), .D(n19668), .Y(n17375) );
  MUX2X1 U10887 ( .B(n19574), .A(msg[22]), .S(n16983), .Y(n17286) );
  AOI22X1 U10888 ( .A(msg[7]), .B(msg[8]), .C(n19619), .D(n19626), .Y(n17210)
         );
  MUX2X1 U10889 ( .B(n19561), .A(msg[27]), .S(n16990), .Y(n17436) );
  AOI22X1 U10890 ( .A(msg[43]), .B(msg[5]), .C(n19632), .D(n19450), .Y(n17270)
         );
  AOI22X1 U10891 ( .A(msg[19]), .B(msg[40]), .C(n19522), .D(n19583), .Y(n19676) );
  INVX1 U10892 ( .A(n19676), .Y(n19677) );
  FAX1 U10893 ( .A(n17291), .B(n17093), .C(n19677), .YS(n17176) );
  FAX1 U10894 ( .A(n17286), .B(n17436), .C(n17176), .YS(n17177) );
  FAX1 U10895 ( .A(n17280), .B(n17463), .C(n17177), .YS(n17467) );
  INVX1 U10896 ( .A(msg[55]), .Y(n17271) );
  MUX2X1 U10897 ( .B(msg[55]), .A(n17271), .S(n19585), .Y(n17178) );
  MUX2X1 U10898 ( .B(n19597), .A(msg[15]), .S(n17178), .Y(n17385) );
  INVX1 U10899 ( .A(msg[58]), .Y(n17204) );
  MUX2X1 U10900 ( .B(msg[58]), .A(n17204), .S(n17213), .Y(n19680) );
  AOI22X1 U10901 ( .A(msg[48]), .B(msg[28]), .C(n19559), .D(n17290), .Y(n17221) );
  MUX2X1 U10902 ( .B(msg[39]), .A(n19525), .S(n19677), .Y(n17247) );
  HAX1 U10903 ( .A(n17038), .B(n17247), .YS(n17179) );
  FAX1 U10904 ( .A(n17385), .B(n19680), .C(n17179), .YS(n17198) );
  MUX2X1 U10905 ( .B(n19651), .A(msg[1]), .S(n17194), .Y(n17180) );
  MUX2X1 U10906 ( .B(n19450), .A(msg[43]), .S(n17180), .Y(n17403) );
  HAX1 U10907 ( .A(n17082), .B(n17288), .YS(n17190) );
  MUX2X1 U10908 ( .B(n19565), .A(msg[25]), .S(n17190), .Y(n17182) );
  MUX2X1 U10909 ( .B(n19609), .A(msg[11]), .S(n17182), .Y(n17442) );
  INVX1 U10910 ( .A(n17379), .Y(n17378) );
  HAX1 U10911 ( .A(n17183), .B(n17378), .YS(n17218) );
  AOI22X1 U10912 ( .A(msg[45]), .B(msg[21]), .C(n19576), .D(n17376), .Y(n17184) );
  MUX2X1 U10913 ( .B(n17185), .A(msg[46]), .S(n17184), .Y(n17186) );
  MUX2X1 U10914 ( .B(msg[49]), .A(n17187), .S(n17186), .Y(n17188) );
  FAX1 U10915 ( .A(n17442), .B(n17218), .C(n17188), .YS(n17189) );
  FAX1 U10916 ( .A(n17198), .B(n17403), .C(n17189), .YS(n17390) );
  NAND3X1 U10917 ( .A(n16904), .B(n17467), .C(n17390), .Y(n18748) );
  MUX2X1 U10918 ( .B(n17199), .A(msg[57]), .S(n17190), .Y(n17459) );
  HAX1 U10919 ( .A(n17192), .B(n16592), .YS(n17414) );
  AOI22X1 U10920 ( .A(msg[31]), .B(msg[9]), .C(n19615), .D(n19551), .Y(n17193)
         );
  FAX1 U10921 ( .A(n17194), .B(n17093), .C(n16593), .YS(n17195) );
  MUX2X1 U10922 ( .B(n19509), .A(msg[41]), .S(n17195), .Y(n17196) );
  FAX1 U10923 ( .A(n17220), .B(n17414), .C(n17196), .YS(n17197) );
  FAX1 U10924 ( .A(n17198), .B(n17459), .C(n17197), .YS(n18323) );
  AOI22X1 U10925 ( .A(msg[57]), .B(msg[26]), .C(n19563), .D(n17199), .Y(n17275) );
  MUX2X1 U10926 ( .B(n19546), .A(msg[32]), .S(msg[50]), .Y(n19679) );
  FAX1 U10927 ( .A(n17200), .B(n17025), .C(n19679), .YS(n17203) );
  AOI22X1 U10928 ( .A(msg[34]), .B(msg[4]), .C(n19637), .D(n19539), .Y(n17233)
         );
  MUX2X1 U10929 ( .B(n17231), .A(msg[56]), .S(n17030), .Y(n17202) );
  HAX1 U10930 ( .A(n17432), .B(n17247), .YS(n17201) );
  FAX1 U10931 ( .A(n17203), .B(n17202), .C(n17201), .YS(n17208) );
  MUX2X1 U10932 ( .B(msg[58]), .A(n17204), .S(n17436), .Y(n17370) );
  INVX1 U10933 ( .A(n17370), .Y(n17205) );
  HAX1 U10934 ( .A(n17081), .B(n17205), .YS(n17206) );
  MUX2X1 U10935 ( .B(n19629), .A(msg[6]), .S(n17206), .Y(n17249) );
  INVX1 U10936 ( .A(n17249), .Y(n17207) );
  FAX1 U10937 ( .A(n17209), .B(n17208), .C(n17207), .YS(n18329) );
  XNOR2X1 U10938 ( .A(n16990), .B(n17418), .Y(n17279) );
  MUX2X1 U10939 ( .B(msg[36]), .A(n19533), .S(n17279), .Y(n17238) );
  MUX2X1 U10940 ( .B(msg[0]), .A(n19656), .S(n17211), .Y(n17212) );
  MUX2X1 U10941 ( .B(n19637), .A(msg[4]), .S(n17212), .Y(n19689) );
  MUX2X1 U10942 ( .B(msg[52]), .A(n17213), .S(n19689), .Y(n17214) );
  FAX1 U10943 ( .A(n17215), .B(n17238), .C(n17214), .YS(n17216) );
  FAX1 U10944 ( .A(n17218), .B(n17217), .C(n17216), .YS(n17219) );
  FAX1 U10945 ( .A(n17038), .B(n17220), .C(n17219), .YS(n18333) );
  NAND2X1 U10946 ( .A(n18329), .B(n18333), .Y(n17600) );
  OR2X1 U10947 ( .A(n18323), .B(n17600), .Y(n17628) );
  INVX1 U10948 ( .A(n17628), .Y(n17597) );
  INVX1 U10949 ( .A(n17467), .Y(n17594) );
  INVX1 U10950 ( .A(n17222), .Y(n17598) );
  INVX1 U10951 ( .A(n17588), .Y(n17602) );
  NAND2X1 U10952 ( .A(n17597), .B(n18322), .Y(n17666) );
  AOI21X1 U10953 ( .A(n17224), .B(n17342), .C(n17002), .Y(n17307) );
  INVX1 U10954 ( .A(\lamb/scale_ds1/genblk1[3].mult/added[3] ), .Y(n17344) );
  OR2X1 U10955 ( .A(n17344), .B(\add_x_71/n1 ), .Y(n17225) );
  AOI22X1 U10956 ( .A(\lamb/scale_ds1/genblk1[3].mult/added[4] ), .B(
        \lamb/scale_ds1/genblk1[3].mult/added[3] ), .C(n17065), .D(n17225), 
        .Y(n17357) );
  AOI21X1 U10957 ( .A(\lamb/scale_ds1/genblk1[3].mult/added[1] ), .B(n16582), 
        .C(\lamb/scale_ds1/genblk1[3].mult/added[2] ), .Y(n17227) );
  NAND3X1 U10958 ( .A(\lamb/scale_ds1/genblk1[3].mult/added[4] ), .B(
        \add_x_71/n1 ), .C(\lamb/scale_ds1/genblk1[3].mult/added[3] ), .Y(
        n17311) );
  OR2X1 U10959 ( .A(\lamb/scale_ds1/genblk1[3].mult/added[4] ), .B(
        \add_x_71/n1 ), .Y(n17312) );
  OR2X1 U10960 ( .A(n17312), .B(\lamb/scale_ds1/genblk1[3].mult/added[3] ), 
        .Y(n17316) );
  NAND2X1 U10961 ( .A(\lamb/scale_ds1/genblk1[3].mult/added[3] ), .B(n17312), 
        .Y(n17308) );
  INVX1 U10962 ( .A(n17308), .Y(n17226) );
  INVX1 U10963 ( .A(\lamb/scale_ds1/genblk1[3].mult/added[1] ), .Y(n17347) );
  NAND3X1 U10964 ( .A(n17226), .B(n17347), .C(n17065), .Y(n17361) );
  AOI22X1 U10965 ( .A(n17227), .B(n16659), .C(n17310), .D(n17361), .Y(n17349)
         );
  OR2X1 U10966 ( .A(\lamb/scale_ds1/genblk1[3].mult/added[1] ), .B(n16659), 
        .Y(n17230) );
  NAND3X1 U10967 ( .A(n16659), .B(\lamb/scale_ds1/genblk1[3].mult/added[2] ), 
        .C(\lamb/scale_ds1/genblk1[3].mult/added[1] ), .Y(n17228) );
  NAND2X1 U10968 ( .A(n17228), .B(n17316), .Y(n17345) );
  INVX1 U10969 ( .A(n17345), .Y(n17229) );
  NAND2X1 U10970 ( .A(n17230), .B(n17229), .Y(n17305) );
  AOI22X1 U10971 ( .A(msg[5]), .B(msg[42]), .C(n19670), .D(n19632), .Y(n17373)
         );
  MUX2X1 U10972 ( .B(n17231), .A(msg[56]), .S(n17411), .Y(n17232) );
  MUX2X1 U10973 ( .B(msg[23]), .A(n19572), .S(n17232), .Y(n17434) );
  FAX1 U10974 ( .A(n17234), .B(n17030), .C(n17434), .YS(n17235) );
  FAX1 U10975 ( .A(n17236), .B(n16716), .C(n17235), .YS(n17237) );
  FAX1 U10976 ( .A(n17463), .B(n17238), .C(n17237), .YS(n18375) );
  INVX1 U10977 ( .A(n18375), .Y(n18381) );
  INVX1 U10978 ( .A(\lamb/scale_ts0/genblk1[2].mult/added[3] ), .Y(n17256) );
  NOR2X1 U10979 ( .A(n17256), .B(n17095), .Y(n17239) );
  INVX1 U10980 ( .A(\lamb/scale_ts0/genblk1[2].mult/added[1] ), .Y(n17263) );
  NAND2X1 U10981 ( .A(\lamb/scale_ts0/genblk1[2].mult/added[4] ), .B(
        \add_x_77/n1 ), .Y(n17255) );
  NAND3X1 U10982 ( .A(n17239), .B(n17263), .C(n17255), .Y(n17258) );
  AOI21X1 U10983 ( .A(\add_x_77/n1 ), .B(
        \lamb/scale_ts0/genblk1[2].mult/added[4] ), .C(
        \lamb/scale_ts0/genblk1[2].mult/added[3] ), .Y(n17241) );
  INVX1 U10984 ( .A(n17241), .Y(n17262) );
  OAI21X1 U10985 ( .A(n17256), .B(n17095), .C(n17262), .Y(n17268) );
  INVX1 U10986 ( .A(n17268), .Y(n17300) );
  OAI21X1 U10987 ( .A(\lamb/scale_ts0/genblk1[2].mult/added[3] ), .B(
        \lamb/scale_ts0/genblk1[2].mult/added[2] ), .C(
        \lamb/scale_ts0/genblk1[2].mult/added[1] ), .Y(n17240) );
  AOI21X1 U10988 ( .A(n17262), .B(n17265), .C(n17240), .Y(n17269) );
  AOI21X1 U10989 ( .A(\lamb/scale_ts0/genblk1[2].mult/added[2] ), .B(n17300), 
        .C(n16922), .Y(n17243) );
  NAND3X1 U10990 ( .A(\lamb/scale_ts0/genblk1[2].mult/added[1] ), .B(n17241), 
        .C(n17264), .Y(n17242) );
  NAND3X1 U10991 ( .A(n17258), .B(n17243), .C(n17242), .Y(n17244) );
  NAND2X1 U10992 ( .A(n18413), .B(n17244), .Y(n17245) );
  HAX1 U10993 ( .A(n18381), .B(n17245), .YS(n19699) );
  MUX2X1 U10994 ( .B(n19527), .A(msg[38]), .S(n17246), .Y(n19674) );
  HAX1 U10995 ( .A(n17247), .B(n17435), .YS(n17272) );
  MUX2X1 U10996 ( .B(n19656), .A(msg[0]), .S(n17248), .Y(n17402) );
  FAX1 U10997 ( .A(n17251), .B(n17250), .C(n17249), .YS(n17252) );
  FAX1 U10998 ( .A(n17272), .B(n17402), .C(n17252), .YS(n17253) );
  FAX1 U10999 ( .A(n17254), .B(n19674), .C(n17253), .YS(n17622) );
  INVX1 U11000 ( .A(n17622), .Y(n18382) );
  AND2X1 U11001 ( .A(n17263), .B(n17262), .Y(n19692) );
  NAND2X1 U11002 ( .A(\lamb/scale_ts0/genblk1[2].mult/added[1] ), .B(
        \lamb/scale_ts0/genblk1[2].mult/added[2] ), .Y(n17257) );
  NAND2X1 U11003 ( .A(n17095), .B(n17256), .Y(n17259) );
  OAI21X1 U11004 ( .A(n17067), .B(n17257), .C(n17259), .Y(n17297) );
  NAND3X1 U11005 ( .A(n17259), .B(n17258), .C(
        \lamb/scale_ts0/genblk1[2].mult/added[2] ), .Y(n17260) );
  OAI21X1 U11006 ( .A(\lamb/scale_ts0/genblk1[2].mult/added[2] ), .B(n17067), 
        .C(n17260), .Y(n17302) );
  OAI21X1 U11007 ( .A(n19692), .B(n17297), .C(n17302), .Y(n19691) );
  NAND2X1 U11008 ( .A(n18413), .B(n19691), .Y(n17261) );
  HAX1 U11009 ( .A(n18382), .B(n17261), .YS(n18336) );
  AOI21X1 U11010 ( .A(n17095), .B(n17263), .C(n17262), .Y(n17266) );
  OAI21X1 U11011 ( .A(n17067), .B(n17266), .C(n17265), .Y(n17267) );
  AOI22X1 U11012 ( .A(\lamb/scale_ts0/genblk1[2].mult/added[1] ), .B(
        \lamb/scale_ts0/genblk1[2].mult/added[2] ), .C(n17268), .D(n17267), 
        .Y(n17298) );
  OAI21X1 U11013 ( .A(n16922), .B(n16366), .C(n18413), .Y(n17282) );
  MUX2X1 U11014 ( .B(msg[45]), .A(n17376), .S(n17093), .Y(n19686) );
  MUX2X1 U11015 ( .B(msg[55]), .A(n17271), .S(n19686), .Y(n17431) );
  HAX1 U11016 ( .A(n17273), .B(n17272), .YS(n17405) );
  MUX2X1 U11017 ( .B(n19529), .A(msg[37]), .S(n17274), .Y(n17277) );
  INVX1 U11018 ( .A(n17025), .Y(n17276) );
  FAX1 U11019 ( .A(msg[35]), .B(n17277), .C(n17276), .YS(n17278) );
  FAX1 U11020 ( .A(n17280), .B(n17279), .C(n17278), .YS(n17281) );
  FAX1 U11021 ( .A(n17431), .B(n17405), .C(n17281), .YS(n18384) );
  INVX1 U11022 ( .A(n18384), .Y(n17642) );
  HAX1 U11023 ( .A(n17282), .B(n17642), .YS(n18337) );
  MUX2X1 U11024 ( .B(msg[53]), .A(n17283), .S(n19686), .Y(n17456) );
  FAX1 U11025 ( .A(n17285), .B(n16714), .C(n17456), .YS(n17421) );
  MUX2X1 U11026 ( .B(n19619), .A(msg[8]), .S(n17286), .Y(n17287) );
  MUX2X1 U11027 ( .B(n19509), .A(msg[41]), .S(n17287), .Y(n17296) );
  MUX2X1 U11028 ( .B(n19605), .A(msg[12]), .S(n17288), .Y(n17289) );
  MUX2X1 U11029 ( .B(n17290), .A(msg[48]), .S(n17289), .Y(n17372) );
  MUX2X1 U11030 ( .B(n19651), .A(msg[1]), .S(n17291), .Y(n17371) );
  HAX1 U11031 ( .A(n17293), .B(n17292), .YS(n17294) );
  FAX1 U11032 ( .A(n17372), .B(n17371), .C(n17294), .YS(n17295) );
  FAX1 U11033 ( .A(n17421), .B(n17296), .C(n17295), .YS(n18380) );
  INVX1 U11034 ( .A(n18380), .Y(n17614) );
  INVX1 U11035 ( .A(n17297), .Y(n17303) );
  AOI22X1 U11036 ( .A(\lamb/scale_ts0/genblk1[2].mult/added[1] ), .B(n17300), 
        .C(n17067), .D(n16366), .Y(n17301) );
  NAND3X1 U11037 ( .A(n17303), .B(n17302), .C(n17301), .Y(n19690) );
  NAND2X1 U11038 ( .A(n16378), .B(n18413), .Y(n17304) );
  HAX1 U11039 ( .A(n17614), .B(n17304), .YS(n18334) );
  NAND2X1 U11040 ( .A(n18336), .B(n17047), .Y(n18342) );
  OAI21X1 U11041 ( .A(n17349), .B(n17305), .C(n17035), .Y(n17306) );
  HAX1 U11042 ( .A(n17307), .B(n17306), .YS(n19703) );
  INVX1 U11043 ( .A(n19703), .Y(n19712) );
  INVX1 U11044 ( .A(\lamb/scale_ds1/genblk1[3].mult/added[2] ), .Y(n17318) );
  NAND2X1 U11045 ( .A(n17318), .B(n17308), .Y(n17309) );
  NAND3X1 U11046 ( .A(\lamb/scale_ds1/genblk1[3].mult/added[1] ), .B(n16899), 
        .C(n17309), .Y(n17359) );
  INVX1 U11047 ( .A(n17359), .Y(n17322) );
  INVX1 U11048 ( .A(n16582), .Y(n17315) );
  NAND2X1 U11049 ( .A(n16659), .B(n17315), .Y(n17314) );
  NAND3X1 U11050 ( .A(n17312), .B(n17344), .C(n17065), .Y(n17313) );
  INVX1 U11051 ( .A(n17313), .Y(n17358) );
  AOI21X1 U11052 ( .A(n17347), .B(n17314), .C(n17358), .Y(n17320) );
  OAI21X1 U11053 ( .A(n17316), .B(n17347), .C(n17315), .Y(n17317) );
  INVX1 U11054 ( .A(n17317), .Y(n17319) );
  AOI22X1 U11055 ( .A(\lamb/scale_ds1/genblk1[3].mult/added[2] ), .B(n16821), 
        .C(n17319), .D(n17318), .Y(n17321) );
  OAI21X1 U11056 ( .A(n17322), .B(n17321), .C(n17035), .Y(n17335) );
  AOI21X1 U11057 ( .A(\lamb/scale_ts1/genblk1[3].mult/added[1] ), .B(
        \lamb/scale_ts1/genblk1[3].mult/added[2] ), .C(n16893), .Y(n17333) );
  AND2X1 U11058 ( .A(n17325), .B(n17324), .Y(n17352) );
  AOI22X1 U11059 ( .A(\lamb/scale_ts1/genblk1[3].mult/added[1] ), .B(n17336), 
        .C(\lamb/scale_ts1/genblk1[3].mult/added[2] ), .D(n17352), .Y(n17331)
         );
  INVX1 U11060 ( .A(\lamb/scale_ts1/genblk1[3].mult/added[2] ), .Y(n17326) );
  NAND2X1 U11061 ( .A(n16476), .B(n17326), .Y(n17328) );
  NAND3X1 U11062 ( .A(n17331), .B(n17330), .C(n17353), .Y(n17332) );
  OAI21X1 U11063 ( .A(n17333), .B(n17332), .C(n17340), .Y(n17334) );
  HAX1 U11064 ( .A(n17335), .B(n17334), .YS(n18155) );
  INVX1 U11065 ( .A(n16422), .Y(n17366) );
  INVX1 U11066 ( .A(n17336), .Y(n17338) );
  OR2X1 U11067 ( .A(\lamb/scale_ts1/genblk1[3].mult/added[1] ), .B(n17352), 
        .Y(n17337) );
  NAND3X1 U11068 ( .A(n17339), .B(n17338), .C(n17337), .Y(n17341) );
  AOI21X1 U11069 ( .A(n17342), .B(n17341), .C(n17002), .Y(n17351) );
  NAND2X1 U11070 ( .A(n17344), .B(n17065), .Y(n17346) );
  AOI21X1 U11071 ( .A(n17347), .B(n17346), .C(n17345), .Y(n17348) );
  OAI21X1 U11072 ( .A(n17349), .B(n17348), .C(n17035), .Y(n17350) );
  HAX1 U11073 ( .A(n17351), .B(n17350), .YS(n19713) );
  INVX1 U11074 ( .A(n19713), .Y(n18122) );
  AOI22X1 U11075 ( .A(\lamb/scale_ts1/genblk1[3].mult/added[1] ), .B(n17352), 
        .C(\lamb/scale_ts1/genblk1[3].mult/added[2] ), .D(n17323), .Y(n17354)
         );
  NAND3X1 U11076 ( .A(n17355), .B(n17354), .C(n17353), .Y(n17356) );
  NAND2X1 U11077 ( .A(n17340), .B(n17356), .Y(n17365) );
  AOI22X1 U11078 ( .A(\lamb/scale_ds1/genblk1[3].mult/added[1] ), .B(n17358), 
        .C(\lamb/scale_ds1/genblk1[3].mult/added[2] ), .D(n16582), .Y(n17360)
         );
  NAND3X1 U11079 ( .A(n17361), .B(n17360), .C(n17359), .Y(n17363) );
  NAND2X1 U11080 ( .A(n17363), .B(n17035), .Y(n17364) );
  HAX1 U11081 ( .A(n17365), .B(n17364), .YS(n19711) );
  INVX1 U11082 ( .A(n19711), .Y(n19772) );
  NAND2X1 U11083 ( .A(n18122), .B(n19703), .Y(n19701) );
  INVX1 U11084 ( .A(n19701), .Y(n19709) );
  NAND2X1 U11085 ( .A(n19711), .B(n18155), .Y(n19714) );
  AOI22X1 U11086 ( .A(n17366), .B(n16897), .C(n19709), .D(n19714), .Y(n17367)
         );
  INVX1 U11087 ( .A(n18155), .Y(n19710) );
  NAND2X1 U11088 ( .A(n19772), .B(n19710), .Y(n17512) );
  AND2X1 U11089 ( .A(n17367), .B(n17512), .Y(
        \lamb/scale_bs2/genblk1[1].mult/added[3] ) );
  INVX1 U11090 ( .A(n17579), .Y(n17595) );
  NAND2X1 U11091 ( .A(n17595), .B(n16642), .Y(n17587) );
  OAI21X1 U11092 ( .A(n17585), .B(n16570), .C(n17587), .Y(n17368) );
  AND2X1 U11093 ( .A(n16548), .B(n17368), .Y(n16314) );
  MUX2X1 U11094 ( .B(msg[13]), .A(n19601), .S(n17370), .Y(n17420) );
  MUX2X1 U11095 ( .B(n19647), .A(msg[2]), .S(n17371), .Y(n17441) );
  MUX2X1 U11096 ( .B(n19576), .A(msg[21]), .S(n17441), .Y(n19696) );
  FAX1 U11097 ( .A(n17039), .B(n16716), .C(n17372), .YS(n17384) );
  MUX2X1 U11098 ( .B(n17376), .A(msg[45]), .S(n16983), .Y(n17377) );
  MUX2X1 U11099 ( .B(n17379), .A(n17378), .S(n17377), .Y(n17380) );
  MUX2X1 U11100 ( .B(n17382), .A(n17381), .S(n17380), .Y(n17383) );
  FAX1 U11101 ( .A(n17385), .B(n17384), .C(n17383), .YS(n17386) );
  FAX1 U11102 ( .A(n17420), .B(n19696), .C(n17386), .YS(n17591) );
  OAI21X1 U11103 ( .A(n17591), .B(n17716), .C(n16485), .Y(
        \lamb/scale_ts0/genblk1[2].mult/logA[0] ) );
  AND2X1 U11104 ( .A(n17630), .B(\lamb/scale_ts0/genblk1[2].mult/logA[0] ), 
        .Y(\lamb/scale_ts1/genblk1[3].mult/logA[0] ) );
  INVX1 U11105 ( .A(n18322), .Y(n17596) );
  INVX1 U11106 ( .A(n18323), .Y(n17599) );
  AOI21X1 U11107 ( .A(n16482), .B(n16982), .C(n18333), .Y(n17387) );
  INVX1 U11108 ( .A(n18329), .Y(n18330) );
  NAND2X1 U11109 ( .A(n17596), .B(n18330), .Y(n18320) );
  INVX1 U11110 ( .A(n18320), .Y(n18327) );
  OR2X1 U11111 ( .A(n17387), .B(n18327), .Y(
        \lamb/scale_ts1/genblk1[0].mult/logB[0] ) );
  AOI21X1 U11112 ( .A(n17589), .B(n17590), .C(n17390), .Y(n17388) );
  MUX2X1 U11113 ( .B(n16485), .A(n17594), .S(n17388), .Y(n18298) );
  AND2X1 U11114 ( .A(n16709), .B(n17630), .Y(
        \lamb/scale_ls2/genblk1[1].mult/logA[2] ) );
  INVX1 U11115 ( .A(n17390), .Y(n17603) );
  OAI21X1 U11116 ( .A(n17716), .B(n16344), .C(n17589), .Y(n17392) );
  AOI22X1 U11117 ( .A(n16344), .B(n17716), .C(n17392), .D(n17467), .Y(
        \lamb/scale_ts0/genblk1[2].mult/logA[1] ) );
  OR2X1 U11118 ( .A(\add_x_78/n1 ), .B(
        \lamb/scale_ts0/genblk1[1].mult/added[4] ), .Y(n17407) );
  NAND2X1 U11119 ( .A(\lamb/scale_ts0/genblk1[1].mult/added[3] ), .B(n17407), 
        .Y(n17427) );
  INVX1 U11120 ( .A(n17427), .Y(n17446) );
  NAND2X1 U11121 ( .A(\add_x_78/n1 ), .B(
        \lamb/scale_ts0/genblk1[1].mult/added[4] ), .Y(n17394) );
  NOR2X1 U11122 ( .A(n17446), .B(n16524), .Y(n17455) );
  OR2X1 U11123 ( .A(n17407), .B(\lamb/scale_ts0/genblk1[1].mult/added[3] ), 
        .Y(n17447) );
  INVX1 U11124 ( .A(\lamb/scale_ts0/genblk1[1].mult/added[1] ), .Y(n17445) );
  NAND3X1 U11125 ( .A(\lamb/scale_ts0/genblk1[1].mult/added[3] ), .B(
        \add_x_78/n1 ), .C(\lamb/scale_ts0/genblk1[1].mult/added[4] ), .Y(
        n17444) );
  INVX1 U11126 ( .A(\lamb/scale_ts0/genblk1[1].mult/added[2] ), .Y(n17426) );
  AOI22X1 U11127 ( .A(n17423), .B(n17430), .C(n16652), .D(n17426), .Y(n17410)
         );
  AOI21X1 U11128 ( .A(n17455), .B(\lamb/scale_ts0/genblk1[1].mult/added[1] ), 
        .C(n17410), .Y(n17397) );
  MUX2X1 U11129 ( .B(n17445), .A(\lamb/scale_ts0/genblk1[1].mult/added[1] ), 
        .S(n16652), .Y(n17395) );
  OAI21X1 U11130 ( .A(n17426), .B(n17395), .C(n17447), .Y(n17408) );
  INVX1 U11131 ( .A(n17408), .Y(n17396) );
  NOR2X1 U11132 ( .A(n18384), .B(n18380), .Y(n18377) );
  NAND2X1 U11133 ( .A(n18384), .B(n18380), .Y(n18374) );
  AOI21X1 U11134 ( .A(n17622), .B(n18374), .C(n18381), .Y(n18378) );
  AOI21X1 U11135 ( .A(n17397), .B(n17396), .C(n16638), .Y(n17406) );
  HAX1 U11136 ( .A(n17399), .B(n16591), .YS(n17416) );
  MUX2X1 U11137 ( .B(msg[2]), .A(n19647), .S(n17416), .Y(n17400) );
  MUX2X1 U11138 ( .B(n19668), .A(msg[59]), .S(n17400), .Y(n17401) );
  FAX1 U11139 ( .A(n17403), .B(n17402), .C(n17401), .YS(n17404) );
  FAX1 U11140 ( .A(n17462), .B(n17405), .C(n17404), .YS(n17499) );
  HAX1 U11141 ( .A(n17406), .B(n17499), .YS(n18348) );
  INVX1 U11142 ( .A(n17630), .Y(n18752) );
  NAND2X1 U11143 ( .A(n18752), .B(n17594), .Y(n17605) );
  AOI22X1 U11144 ( .A(n18380), .B(n17738), .C(n18348), .D(n17123), .Y(n18216)
         );
  NAND2X1 U11145 ( .A(n18752), .B(n17603), .Y(n18302) );
  OAI21X1 U11146 ( .A(n18752), .B(n18382), .C(n18302), .Y(n17665) );
  AOI21X1 U11147 ( .A(n17445), .B(n17019), .C(n17408), .Y(n17409) );
  OAI21X1 U11148 ( .A(n17410), .B(n17409), .C(n17451), .Y(n17422) );
  AOI22X1 U11149 ( .A(msg[25]), .B(msg[28]), .C(n19559), .D(n19565), .Y(n17415) );
  HAX1 U11150 ( .A(n17412), .B(n17411), .YS(n17413) );
  FAX1 U11151 ( .A(n16712), .B(n17414), .C(n17413), .YS(n17417) );
  FAX1 U11152 ( .A(n17418), .B(n17417), .C(n17416), .YS(n17419) );
  FAX1 U11153 ( .A(n17421), .B(n17420), .C(n17419), .YS(n17502) );
  HAX1 U11154 ( .A(n17422), .B(n17502), .YS(n18346) );
  AOI22X1 U11155 ( .A(n18156), .B(n17665), .C(n18346), .D(n17123), .Y(n18212)
         );
  INVX1 U11156 ( .A(n16663), .Y(n18217) );
  OR2X1 U11157 ( .A(n16750), .B(n18217), .Y(n18221) );
  AND2X1 U11158 ( .A(n18752), .B(n17590), .Y(n18296) );
  AOI21X1 U11159 ( .A(n17630), .B(n18381), .C(n18296), .Y(n19756) );
  INVX1 U11160 ( .A(n17079), .Y(n18307) );
  OAI21X1 U11161 ( .A(n17446), .B(\lamb/scale_ts0/genblk1[1].mult/added[2] ), 
        .C(n16882), .Y(n17424) );
  NAND2X1 U11162 ( .A(n17019), .B(n17424), .Y(n17428) );
  AOI22X1 U11163 ( .A(\lamb/scale_ts0/genblk1[1].mult/added[1] ), .B(n17428), 
        .C(n16327), .D(n17427), .Y(n17429) );
  AOI21X1 U11164 ( .A(n17430), .B(n17429), .C(n16638), .Y(n17443) );
  FAX1 U11165 ( .A(n17433), .B(n17432), .C(n17431), .YS(n17438) );
  FAX1 U11166 ( .A(n17436), .B(n17435), .C(n17434), .YS(n17437) );
  FAX1 U11167 ( .A(n17439), .B(n17438), .C(n17437), .YS(n17440) );
  FAX1 U11168 ( .A(n17442), .B(n17441), .C(n17440), .YS(n17503) );
  INVX1 U11169 ( .A(n17503), .Y(n17631) );
  HAX1 U11170 ( .A(n17443), .B(n17631), .YS(n18344) );
  AOI22X1 U11171 ( .A(n18156), .B(n18307), .C(n18344), .D(n17123), .Y(n18224)
         );
  AOI21X1 U11172 ( .A(n18221), .B(n16601), .C(n16761), .Y(n17465) );
  NAND2X1 U11173 ( .A(n18752), .B(n17589), .Y(n18300) );
  OAI21X1 U11174 ( .A(n18752), .B(n17642), .C(n18300), .Y(n19753) );
  AND2X1 U11175 ( .A(n17445), .B(n16652), .Y(n17450) );
  AOI21X1 U11176 ( .A(\lamb/scale_ts0/genblk1[1].mult/added[1] ), .B(n17446), 
        .C(\lamb/scale_ts0/genblk1[1].mult/added[2] ), .Y(n17448) );
  AOI22X1 U11177 ( .A(n17450), .B(n17019), .C(n17448), .D(n17447), .Y(n17454)
         );
  AOI21X1 U11178 ( .A(\lamb/scale_ts0/genblk1[1].mult/added[1] ), .B(n16327), 
        .C(n16638), .Y(n17453) );
  OAI21X1 U11179 ( .A(n17455), .B(n17454), .C(n17453), .Y(n17464) );
  MUX2X1 U11180 ( .B(n17457), .A(msg[51]), .S(n17456), .Y(n17458) );
  FAX1 U11181 ( .A(n17081), .B(n17459), .C(n17458), .YS(n17461) );
  FAX1 U11182 ( .A(n17463), .B(n17462), .C(n17461), .YS(n17498) );
  INVX1 U11183 ( .A(n17498), .Y(n17643) );
  HAX1 U11184 ( .A(n17464), .B(n17643), .YS(n19719) );
  AOI22X1 U11185 ( .A(n18156), .B(n19753), .C(n19719), .D(n17123), .Y(n18222)
         );
  OR2X1 U11186 ( .A(n17465), .B(n16650), .Y(n9906) );
  HAX1 U11187 ( .A(n17643), .B(n16978), .YS(n17466) );
  INVX1 U11188 ( .A(n17502), .Y(n17621) );
  INVX1 U11189 ( .A(n17499), .Y(n17615) );
  OAI21X1 U11190 ( .A(n17503), .B(n17466), .C(n16386), .Y(
        \lamb/scale_ts0/genblk1[0].mult/logA[3] ) );
  INVX1 U11191 ( .A(\lamb/scale_ts0/genblk1[0].mult/logA[3] ), .Y(n17468) );
  NAND3X1 U11192 ( .A(n17468), .B(n17615), .C(n17643), .Y(n18749) );
  INVX1 U11193 ( .A(n16479), .Y(n18278) );
  NOR2X1 U11194 ( .A(\lamb/scale_ts1/genblk1[0].mult/added[4] ), .B(
        \add_x_70/n1 ), .Y(n17474) );
  INVX1 U11195 ( .A(n17474), .Y(n17471) );
  AOI21X1 U11196 ( .A(\add_x_70/n1 ), .B(
        \lamb/scale_ts1/genblk1[0].mult/added[4] ), .C(
        \lamb/scale_ts1/genblk1[0].mult/added[3] ), .Y(n17469) );
  AOI21X1 U11197 ( .A(\lamb/scale_ts1/genblk1[0].mult/added[3] ), .B(n17471), 
        .C(n17469), .Y(n17490) );
  NAND3X1 U11198 ( .A(\lamb/scale_ts1/genblk1[0].mult/added[4] ), .B(
        \add_x_70/n1 ), .C(\lamb/scale_ts1/genblk1[0].mult/added[3] ), .Y(
        n17470) );
  INVX1 U11199 ( .A(n17470), .Y(n17482) );
  OR2X1 U11200 ( .A(\lamb/scale_ts1/genblk1[0].mult/added[2] ), .B(n17482), 
        .Y(n17481) );
  OR2X1 U11201 ( .A(n17471), .B(\lamb/scale_ts1/genblk1[0].mult/added[3] ), 
        .Y(n17485) );
  NAND3X1 U11202 ( .A(\lamb/scale_ts1/genblk1[0].mult/added[3] ), .B(n17471), 
        .C(n16628), .Y(n17492) );
  AOI21X1 U11203 ( .A(\lamb/scale_ts1/genblk1[0].mult/added[4] ), .B(
        \add_x_70/n1 ), .C(n16603), .Y(n17475) );
  AOI21X1 U11204 ( .A(n17481), .B(n16817), .C(n17475), .Y(n17486) );
  AND2X1 U11205 ( .A(\lamb/scale_ts1/genblk1[0].mult/added[4] ), .B(
        \add_x_70/n1 ), .Y(n17473) );
  NOR3X1 U11206 ( .A(n17474), .B(\lamb/scale_ts1/genblk1[0].mult/added[3] ), 
        .C(n17473), .Y(n17488) );
  INVX1 U11207 ( .A(n17488), .Y(n17478) );
  INVX1 U11208 ( .A(\lamb/scale_ts1/genblk1[0].mult/added[1] ), .Y(n17477) );
  INVX1 U11209 ( .A(n17475), .Y(n17476) );
  AOI22X1 U11210 ( .A(n16452), .B(n17478), .C(n17477), .D(n17476), .Y(n17479)
         );
  AOI21X1 U11211 ( .A(\lamb/scale_ts1/genblk1[0].mult/added[2] ), .B(n16613), 
        .C(n17479), .Y(n18275) );
  INVX1 U11212 ( .A(n18275), .Y(n18287) );
  INVX1 U11213 ( .A(n16452), .Y(n17480) );
  OAI21X1 U11214 ( .A(n16628), .B(n17482), .C(n17485), .Y(n18286) );
  NAND3X1 U11215 ( .A(n18287), .B(n17016), .C(n18286), .Y(n18282) );
  INVX1 U11216 ( .A(n18286), .Y(n17483) );
  AOI21X1 U11217 ( .A(\lamb/scale_ts1/genblk1[0].mult/added[1] ), .B(n17483), 
        .C(n17488), .Y(n18268) );
  NAND2X1 U11218 ( .A(n17016), .B(n17483), .Y(n17484) );
  AOI21X1 U11219 ( .A(\lamb/scale_ts1/genblk1[0].mult/added[1] ), .B(n16613), 
        .C(n17484), .Y(n18273) );
  OR2X1 U11220 ( .A(n16603), .B(n16609), .Y(n17487) );
  NAND2X1 U11221 ( .A(n18273), .B(n17487), .Y(n17495) );
  AOI22X1 U11222 ( .A(n16613), .B(n16628), .C(
        \lamb/scale_ts1/genblk1[0].mult/added[2] ), .D(n17488), .Y(n17491) );
  OAI21X1 U11223 ( .A(n16603), .B(n16609), .C(n17491), .Y(n17493) );
  AOI21X1 U11224 ( .A(\lamb/scale_ts1/genblk1[0].mult/added[1] ), .B(n16609), 
        .C(n17493), .Y(n18288) );
  INVX1 U11225 ( .A(n17075), .Y(n18284) );
  NAND2X1 U11226 ( .A(n18284), .B(n17495), .Y(n18269) );
  NAND3X1 U11227 ( .A(n18282), .B(n16968), .C(n18269), .Y(n17496) );
  AND2X1 U11228 ( .A(n18278), .B(n17496), .Y(
        \lamb/scale_ds2/genblk1[1].mult/logA[0] ) );
  OAI21X1 U11229 ( .A(n17503), .B(n17500), .C(n16605), .Y(
        \lamb/scale_ts0/genblk1[0].mult/logA[0] ) );
  AND2X1 U11230 ( .A(n18752), .B(\lamb/scale_ts0/genblk1[0].mult/logA[0] ), 
        .Y(\lamb/scale_ts1/genblk1[0].mult/logA[0] ) );
  AND2X1 U11231 ( .A(n18752), .B(\lamb/scale_ts0/genblk1[0].mult/logA[3] ), 
        .Y(\lamb/scale_ts1/genblk1[0].mult/logA[3] ) );
  NOR2X1 U11232 ( .A(n17502), .B(n17631), .Y(n17505) );
  NAND3X1 U11233 ( .A(n17621), .B(n17503), .C(n16605), .Y(n17507) );
  OAI21X1 U11234 ( .A(n17505), .B(n16605), .C(n17507), .Y(n17506) );
  AOI21X1 U11235 ( .A(n17643), .B(n16328), .C(n17506), .Y(
        \lamb/scale_ts0/genblk1[0].mult/logA[2] ) );
  AND2X1 U11236 ( .A(n18752), .B(n16710), .Y(
        \lamb/scale_ts1/genblk1[0].mult/logA[2] ) );
  AOI22X1 U11237 ( .A(n17615), .B(n17643), .C(n16328), .D(n17507), .Y(
        \lamb/scale_ts0/genblk1[0].mult/logA[1] ) );
  INVX1 U11238 ( .A(\lamb/scale_ls2/genblk1[0].mult/added[1] ), .Y(n17563) );
  OR2X1 U11239 ( .A(\lamb/scale_ls2/genblk1[0].mult/added[4] ), .B(
        \add_x_66/n1 ), .Y(n17531) );
  INVX1 U11240 ( .A(n17531), .Y(n17509) );
  AOI21X1 U11241 ( .A(\add_x_66/n1 ), .B(
        \lamb/scale_ls2/genblk1[0].mult/added[4] ), .C(n17509), .Y(n17542) );
  AND2X1 U11242 ( .A(n17563), .B(n16636), .Y(n17545) );
  INVX1 U11243 ( .A(\lamb/scale_ls2/genblk1[0].mult/added[2] ), .Y(n17532) );
  NAND2X1 U11244 ( .A(\lamb/scale_ls2/genblk1[0].mult/added[3] ), .B(n17532), 
        .Y(n17564) );
  NOR3X1 U11245 ( .A(\lamb/scale_ls2/genblk1[0].mult/added[3] ), .B(
        \lamb/scale_ls2/genblk1[0].mult/added[4] ), .C(\add_x_66/n1 ), .Y(
        n17561) );
  NAND3X1 U11246 ( .A(\lamb/scale_ls2/genblk1[0].mult/added[3] ), .B(
        \lamb/scale_ls2/genblk1[0].mult/added[4] ), .C(\add_x_66/n1 ), .Y(
        n17533) );
  AOI22X1 U11247 ( .A(n17545), .B(n17564), .C(n16960), .D(n16343), .Y(n17511)
         );
  INVX1 U11248 ( .A(n17561), .Y(n17510) );
  OAI21X1 U11249 ( .A(n17052), .B(\lamb/scale_ls2/genblk1[0].mult/added[2] ), 
        .C(n17510), .Y(n17540) );
  NAND2X1 U11250 ( .A(n17052), .B(n17532), .Y(n17560) );
  NAND2X1 U11251 ( .A(n17540), .B(n17560), .Y(n17543) );
  NAND2X1 U11252 ( .A(n17511), .B(n17543), .Y(n17520) );
  OR2X1 U11253 ( .A(n18122), .B(n17512), .Y(n17608) );
  INVX1 U11254 ( .A(n17608), .Y(n17609) );
  NAND2X1 U11255 ( .A(n17630), .B(n16619), .Y(n17538) );
  INVX1 U11256 ( .A(n17538), .Y(n17572) );
  NOR2X1 U11257 ( .A(\lamb/scale_bs2/genblk1[0].mult/added[4] ), .B(
        \add_x_63/n1 ), .Y(n17515) );
  INVX1 U11258 ( .A(\lamb/scale_bs2/genblk1[0].mult/added[3] ), .Y(n17513) );
  NAND3X1 U11259 ( .A(\lamb/scale_bs2/genblk1[0].mult/added[3] ), .B(
        \lamb/scale_bs2/genblk1[0].mult/added[4] ), .C(\add_x_63/n1 ), .Y(
        n17570) );
  INVX1 U11260 ( .A(n16741), .Y(n17525) );
  AOI22X1 U11261 ( .A(n17522), .B(\lamb/scale_bs2/genblk1[0].mult/added[2] ), 
        .C(n17525), .D(\lamb/scale_bs2/genblk1[0].mult/added[1] ), .Y(n17518)
         );
  INVX1 U11262 ( .A(\lamb/scale_bs2/genblk1[0].mult/added[2] ), .Y(n17571) );
  INVX1 U11263 ( .A(\lamb/scale_bs2/genblk1[0].mult/added[1] ), .Y(n17550) );
  NAND2X1 U11264 ( .A(n16741), .B(n17550), .Y(n17514) );
  NAND3X1 U11265 ( .A(n17036), .B(n17571), .C(n17514), .Y(n17517) );
  AOI21X1 U11266 ( .A(\add_x_63/n1 ), .B(
        \lamb/scale_bs2/genblk1[0].mult/added[4] ), .C(n17515), .Y(n17521) );
  NAND3X1 U11267 ( .A(n16521), .B(n17550), .C(n16962), .Y(n17516) );
  NAND3X1 U11268 ( .A(n17518), .B(n17517), .C(n17516), .Y(n17519) );
  AOI22X1 U11269 ( .A(n18303), .B(n17520), .C(n17572), .D(n17519), .Y(n18183)
         );
  NAND2X1 U11270 ( .A(\lamb/scale_bs2/genblk1[0].mult/added[3] ), .B(n16521), 
        .Y(n17549) );
  MUX2X1 U11271 ( .B(\lamb/scale_bs2/genblk1[0].mult/added[2] ), .A(
        \lamb/scale_bs2/genblk1[0].mult/added[1] ), .S(n16467), .Y(n17523) );
  NAND2X1 U11272 ( .A(n16431), .B(n17036), .Y(n17548) );
  AOI22X1 U11273 ( .A(\lamb/scale_bs2/genblk1[0].mult/added[2] ), .B(
        \lamb/scale_bs2/genblk1[0].mult/added[1] ), .C(n17523), .D(n17548), 
        .Y(n17574) );
  AOI21X1 U11274 ( .A(n17525), .B(n17524), .C(n16431), .Y(n17527) );
  NAND2X1 U11275 ( .A(n16741), .B(\lamb/scale_bs2/genblk1[0].mult/added[2] ), 
        .Y(n17526) );
  AOI22X1 U11276 ( .A(n16741), .B(n17550), .C(n16838), .D(n17526), .Y(n17528)
         );
  AOI21X1 U11277 ( .A(n16962), .B(n16467), .C(n17528), .Y(n17539) );
  NAND3X1 U11278 ( .A(\lamb/scale_ls2/genblk1[0].mult/added[3] ), .B(
        \lamb/scale_ls2/genblk1[0].mult/added[2] ), .C(n17531), .Y(n17535) );
  NAND2X1 U11279 ( .A(n16636), .B(n17532), .Y(n17568) );
  NAND3X1 U11280 ( .A(n17568), .B(n17052), .C(
        \lamb/scale_ls2/genblk1[0].mult/added[1] ), .Y(n17534) );
  OAI21X1 U11281 ( .A(\lamb/scale_ls2/genblk1[0].mult/added[1] ), .B(n17535), 
        .C(n17534), .Y(n17536) );
  OAI21X1 U11282 ( .A(n17540), .B(n17536), .C(n18303), .Y(n17537) );
  OAI21X1 U11283 ( .A(n17539), .B(n17538), .C(n17537), .Y(n18190) );
  INVX1 U11284 ( .A(n16647), .Y(n18187) );
  INVX1 U11285 ( .A(n18190), .Y(n18186) );
  OR2X1 U11286 ( .A(n17540), .B(n16636), .Y(n17562) );
  NAND2X1 U11287 ( .A(\lamb/scale_ls2/genblk1[0].mult/added[3] ), .B(
        \lamb/scale_ls2/genblk1[0].mult/added[2] ), .Y(n17541) );
  NAND2X1 U11288 ( .A(n17543), .B(n16894), .Y(n17544) );
  AOI22X1 U11289 ( .A(\lamb/scale_ls2/genblk1[0].mult/added[3] ), .B(n17545), 
        .C(\lamb/scale_ls2/genblk1[0].mult/added[1] ), .D(n17544), .Y(n17546)
         );
  OAI21X1 U11290 ( .A(n16343), .B(n17562), .C(n17546), .Y(n17558) );
  INVX1 U11291 ( .A(n17548), .Y(n17552) );
  INVX1 U11292 ( .A(n17549), .Y(n17551) );
  AOI22X1 U11293 ( .A(\lamb/scale_bs2/genblk1[0].mult/added[2] ), .B(n17552), 
        .C(n17551), .D(n17550), .Y(n17556) );
  OAI21X1 U11294 ( .A(\add_x_63/n1 ), .B(n17571), .C(n16431), .Y(n17555) );
  NAND2X1 U11295 ( .A(\lamb/scale_bs2/genblk1[0].mult/added[3] ), .B(
        \lamb/scale_bs2/genblk1[0].mult/added[2] ), .Y(n17554) );
  NAND3X1 U11296 ( .A(\lamb/scale_bs2/genblk1[0].mult/added[1] ), .B(n17555), 
        .C(n17554), .Y(n17569) );
  NAND2X1 U11297 ( .A(n17556), .B(n17569), .Y(n17557) );
  AOI22X1 U11298 ( .A(n18303), .B(n17558), .C(n17572), .D(n17557), .Y(n18197)
         );
  AOI21X1 U11299 ( .A(n16639), .B(n16380), .C(n17102), .Y(n17577) );
  OAI21X1 U11300 ( .A(n17561), .B(n17560), .C(n16894), .Y(n17567) );
  AOI22X1 U11301 ( .A(n16960), .B(n17564), .C(n17563), .D(n17562), .Y(n17566)
         );
  AOI21X1 U11302 ( .A(n17568), .B(n17567), .C(n17566), .Y(n17576) );
  AOI21X1 U11303 ( .A(n17571), .B(n16741), .C(n17569), .Y(n17573) );
  OAI21X1 U11304 ( .A(n17574), .B(n17573), .C(n17572), .Y(n17575) );
  OAI21X1 U11305 ( .A(n17576), .B(n16661), .C(n17575), .Y(n18194) );
  INVX1 U11306 ( .A(n18194), .Y(n18434) );
  OR2X1 U11307 ( .A(n17577), .B(n16610), .Y(n16300) );
  AND2X1 U11308 ( .A(n18303), .B(\lamb/scale_ts0/genblk1[2].mult/logA[0] ), 
        .Y(\lamb/scale_ls2/genblk1[0].mult/logA[0] ) );
  INVX1 U11309 ( .A(n17578), .Y(n17601) );
  OAI21X1 U11310 ( .A(n17580), .B(n17579), .C(n16622), .Y(n16316) );
  AND2X1 U11311 ( .A(n17628), .B(n16316), .Y(
        \lamb/scale_bs2/genblk1[0].mult/logA[0] ) );
  AND2X1 U11312 ( .A(n16314), .B(n17628), .Y(n16315) );
  OAI21X1 U11313 ( .A(n17588), .B(n17581), .C(n17595), .Y(n17583) );
  AOI22X1 U11314 ( .A(n17581), .B(n17588), .C(n17583), .D(n16642), .Y(
        \lamb/scale_ls1/genblk1[1].mult/added[3] ) );
  AND2X1 U11315 ( .A(n16781), .B(n17628), .Y(
        \lamb/scale_bs2/genblk1[0].mult/logA[3] ) );
  MUX2X1 U11316 ( .B(n17598), .A(n16622), .S(n16570), .Y(n17586) );
  AOI21X1 U11317 ( .A(n17588), .B(n17587), .C(n17586), .Y(
        \lamb/scale_ls1/genblk1[1].mult/added[2] ) );
  AOI21X1 U11318 ( .A(n17589), .B(n17590), .C(n17603), .Y(n17593) );
  NAND2X1 U11319 ( .A(n17590), .B(n17739), .Y(n17592) );
  AOI22X1 U11320 ( .A(n17594), .B(n17593), .C(n17592), .D(n17591), .Y(
        \lamb/scale_ts0/genblk1[2].mult/logA[3] ) );
  INVX1 U11321 ( .A(\lamb/scale_ts0/genblk1[2].mult/logA[3] ), .Y(n18301) );
  OAI21X1 U11322 ( .A(n17608), .B(n16661), .C(n16619), .Y(n18412) );
  INVX1 U11323 ( .A(n18412), .Y(n18414) );
  AND2X1 U11324 ( .A(n18414), .B(\lamb/scale_ls2/genblk1[1].mult/logA[2] ), 
        .Y(\lamb/scale_bs3/genblk1[0].mult/logA[2] ) );
  AND2X1 U11325 ( .A(n18414), .B(\lamb/scale_ts1/genblk1[3].mult/logA[1] ), 
        .Y(\lamb/scale_bs3/genblk1[0].mult/logA[1] ) );
  AND2X1 U11326 ( .A(n18414), .B(\lamb/scale_ts1/genblk1[3].mult/logA[0] ), 
        .Y(\lamb/scale_bs3/genblk1[0].mult/logA[0] ) );
  AND2X1 U11327 ( .A(n18414), .B(n16316), .Y(
        \lamb/scale_bs3/genblk1[1].mult/logA[0] ) );
  AND2X1 U11328 ( .A(n18414), .B(n16781), .Y(
        \lamb/scale_bs3/genblk1[1].mult/logA[3] ) );
  AND2X1 U11329 ( .A(n18414), .B(n16314), .Y(n16303) );
  INVX1 U11330 ( .A(n18333), .Y(n18319) );
  AOI21X1 U11331 ( .A(n17595), .B(n17597), .C(n18319), .Y(n19727) );
  AOI22X1 U11332 ( .A(n17598), .B(n17597), .C(n17596), .D(n16664), .Y(n19731)
         );
  OAI21X1 U11333 ( .A(n17601), .B(n17600), .C(n17599), .Y(n19726) );
  NAND2X1 U11334 ( .A(n16734), .B(n19726), .Y(n19657) );
  NAND3X1 U11335 ( .A(n17603), .B(n17602), .C(n18333), .Y(n17695) );
  INVX1 U11336 ( .A(n16381), .Y(n19730) );
  OR2X1 U11337 ( .A(n16734), .B(n19730), .Y(n19725) );
  OAI21X1 U11338 ( .A(n16745), .B(n16831), .C(n19725), .Y(
        \lamb/scale_ls2/genblk1[0].mult/logB[0] ) );
  OAI21X1 U11339 ( .A(n18752), .B(n17614), .C(n17605), .Y(n17606) );
  INVX1 U11340 ( .A(n17606), .Y(n18309) );
  OR2X1 U11341 ( .A(n17665), .B(n18309), .Y(n19751) );
  AND2X1 U11342 ( .A(n16653), .B(n19751), .Y(n17607) );
  NAND2X1 U11343 ( .A(n19753), .B(n17606), .Y(n17664) );
  OAI21X1 U11344 ( .A(n17079), .B(n17607), .C(n17664), .Y(
        \lamb/scale_ts1/genblk1[2].mult/logA[0] ) );
  AOI21X1 U11345 ( .A(n18412), .B(n16381), .C(n18155), .Y(n18181) );
  AOI22X1 U11346 ( .A(n17609), .B(n16734), .C(n19703), .D(n17608), .Y(n18180)
         );
  INVX1 U11347 ( .A(n16623), .Y(n17612) );
  AOI21X1 U11348 ( .A(n18412), .B(n19726), .C(n18122), .Y(n18179) );
  INVX1 U11349 ( .A(n18179), .Y(n18175) );
  OAI21X1 U11350 ( .A(n18414), .B(n16745), .C(n19772), .Y(n17610) );
  NAND2X1 U11351 ( .A(n16404), .B(n17610), .Y(n18178) );
  INVX1 U11352 ( .A(n17610), .Y(n19770) );
  AOI21X1 U11353 ( .A(n18380), .B(n18382), .C(n17026), .Y(n18376) );
  AOI22X1 U11354 ( .A(n18376), .B(n16340), .C(n16839), .D(n16353), .Y(
        \lamb/scale_ts0/genblk1[1].mult/logA[3] ) );
  MUX2X1 U11355 ( .B(n17615), .A(n17614), .S(n18752), .Y(n19746) );
  INVX1 U11356 ( .A(n16383), .Y(n18369) );
  AND2X1 U11357 ( .A(\lamb/scale_ts0/genblk1[0].mult/added[4] ), .B(
        \add_x_79/n1 ), .Y(n17618) );
  INVX1 U11358 ( .A(n16443), .Y(n17616) );
  OR2X1 U11359 ( .A(\lamb/scale_ts0/genblk1[0].mult/added[4] ), .B(
        \add_x_79/n1 ), .Y(n17623) );
  INVX1 U11360 ( .A(n16488), .Y(n17632) );
  NAND3X1 U11361 ( .A(\lamb/scale_ts0/genblk1[0].mult/added[3] ), .B(
        \lamb/scale_ts0/genblk1[0].mult/added[4] ), .C(\add_x_79/n1 ), .Y(
        n17645) );
  NAND2X1 U11362 ( .A(\lamb/scale_ts0/genblk1[0].mult/added[2] ), .B(
        \lamb/scale_ts0/genblk1[0].mult/added[1] ), .Y(n17638) );
  INVX1 U11363 ( .A(n17638), .Y(n17652) );
  NOR3X1 U11364 ( .A(\lamb/scale_ts0/genblk1[0].mult/added[3] ), .B(
        \lamb/scale_ts0/genblk1[0].mult/added[4] ), .C(\add_x_79/n1 ), .Y(
        n17646) );
  OAI21X1 U11365 ( .A(n17652), .B(n17646), .C(n16627), .Y(n17624) );
  OAI21X1 U11366 ( .A(n16627), .B(\lamb/scale_ts0/genblk1[0].mult/added[1] ), 
        .C(n17624), .Y(n17617) );
  AOI21X1 U11367 ( .A(\lamb/scale_ts0/genblk1[0].mult/added[1] ), .B(n17632), 
        .C(n17617), .Y(n18371) );
  NOR3X1 U11368 ( .A(n17618), .B(\lamb/scale_ts0/genblk1[0].mult/added[1] ), 
        .C(n16611), .Y(n17633) );
  INVX1 U11369 ( .A(n16627), .Y(n17619) );
  INVX1 U11370 ( .A(\lamb/scale_ts0/genblk1[0].mult/added[2] ), .Y(n17636) );
  AOI22X1 U11371 ( .A(\lamb/scale_ts0/genblk1[0].mult/added[2] ), .B(n17633), 
        .C(n17619), .D(n17636), .Y(n17627) );
  NAND2X1 U11372 ( .A(n18369), .B(n16398), .Y(n18355) );
  INVX1 U11373 ( .A(n18355), .Y(n18353) );
  AOI22X1 U11374 ( .A(n19746), .B(n18156), .C(n18353), .D(n17628), .Y(n17620)
         );
  INVX1 U11375 ( .A(n17620), .Y(n18234) );
  MUX2X1 U11376 ( .B(n17622), .A(n17621), .S(n17630), .Y(n18314) );
  AOI22X1 U11377 ( .A(\lamb/scale_ts0/genblk1[0].mult/added[2] ), .B(n17646), 
        .C(\lamb/scale_ts0/genblk1[0].mult/added[1] ), .D(n17624), .Y(n17625)
         );
  OAI21X1 U11378 ( .A(n17652), .B(n17003), .C(n17625), .Y(n18361) );
  INVX1 U11379 ( .A(n18361), .Y(n17626) );
  NAND3X1 U11380 ( .A(n18369), .B(n17628), .C(n17040), .Y(n17629) );
  OAI21X1 U11381 ( .A(n18314), .B(n17123), .C(n17629), .Y(n18228) );
  INVX1 U11382 ( .A(n18228), .Y(n18233) );
  MUX2X1 U11383 ( .B(n18381), .A(n17631), .S(n17630), .Y(n19743) );
  AOI22X1 U11384 ( .A(\lamb/scale_ts0/genblk1[0].mult/added[1] ), .B(n17644), 
        .C(n17652), .D(n17632), .Y(n17641) );
  INVX1 U11385 ( .A(n17633), .Y(n17640) );
  INVX1 U11386 ( .A(\lamb/scale_ts0/genblk1[0].mult/added[1] ), .Y(n17634) );
  AOI22X1 U11387 ( .A(n17636), .B(n16611), .C(n17634), .D(n16488), .Y(n17637)
         );
  OAI21X1 U11388 ( .A(n16443), .B(n17638), .C(n17637), .Y(n17650) );
  NAND3X1 U11389 ( .A(n17641), .B(n17640), .C(n17650), .Y(n18352) );
  AOI22X1 U11390 ( .A(n18156), .B(n19743), .C(n16702), .D(n17123), .Y(n18235)
         );
  MUX2X1 U11391 ( .B(n17643), .A(n17642), .S(n18752), .Y(n19740) );
  NAND2X1 U11392 ( .A(n16627), .B(n17003), .Y(n17647) );
  AOI22X1 U11393 ( .A(\lamb/scale_ts0/genblk1[0].mult/added[2] ), .B(n17647), 
        .C(\lamb/scale_ts0/genblk1[0].mult/added[1] ), .D(n17646), .Y(n17649)
         );
  AND2X1 U11394 ( .A(n17649), .B(n16488), .Y(n17651) );
  OAI21X1 U11395 ( .A(n17652), .B(n17651), .C(n17650), .Y(n18360) );
  AND2X1 U11396 ( .A(n18369), .B(n18360), .Y(n18364) );
  AOI22X1 U11397 ( .A(n18156), .B(n19740), .C(n18364), .D(n17123), .Y(n18236)
         );
  INVX1 U11398 ( .A(n16401), .Y(n18226) );
  NOR2X1 U11399 ( .A(n18234), .B(n18226), .Y(n17950) );
  AOI21X1 U11400 ( .A(n18228), .B(n16574), .C(n16732), .Y(n17949) );
  AOI21X1 U11401 ( .A(n17024), .B(n16732), .C(n17653), .Y(
        \lamb/scale_ts2/genblk1[1].mult/logA[1] ) );
  INVX1 U11402 ( .A(\lamb/scale_ts1/genblk1[2].mult/added[3] ), .Y(n17654) );
  INVX1 U11403 ( .A(n16518), .Y(n17656) );
  NAND2X1 U11404 ( .A(n17015), .B(n17656), .Y(n17698) );
  INVX1 U11405 ( .A(n17698), .Y(n17686) );
  INVX1 U11406 ( .A(n16509), .Y(n17660) );
  NAND2X1 U11407 ( .A(\lamb/scale_ts1/genblk1[2].mult/added[1] ), .B(
        \lamb/scale_ts1/genblk1[2].mult/added[2] ), .Y(n17685) );
  OAI21X1 U11408 ( .A(n17660), .B(n17685), .C(n16320), .Y(n17655) );
  AOI21X1 U11409 ( .A(\lamb/scale_ts1/genblk1[2].mult/added[1] ), .B(n17686), 
        .C(n17655), .Y(n17687) );
  NAND2X1 U11410 ( .A(\lamb/scale_ts1/genblk1[2].mult/added[2] ), .B(n16320), 
        .Y(n17658) );
  INVX1 U11411 ( .A(\lamb/scale_ts1/genblk1[2].mult/added[1] ), .Y(n17689) );
  NAND3X1 U11412 ( .A(n17689), .B(\lamb/scale_ts1/genblk1[2].mult/added[2] ), 
        .C(n17660), .Y(n17657) );
  AOI21X1 U11413 ( .A(n16941), .B(n17657), .C(n17656), .Y(n17729) );
  INVX1 U11414 ( .A(n17658), .Y(n17663) );
  NAND3X1 U11415 ( .A(n16518), .B(n17689), .C(n16509), .Y(n17696) );
  INVX1 U11416 ( .A(\lamb/scale_ts1/genblk1[2].mult/added[2] ), .Y(n17662) );
  NAND2X1 U11417 ( .A(\lamb/scale_ts1/genblk1[2].mult/added[3] ), .B(n17660), 
        .Y(n17661) );
  AOI22X1 U11418 ( .A(n17663), .B(n16364), .C(n17662), .D(n17661), .Y(n17691)
         );
  AOI21X1 U11419 ( .A(n17729), .B(\lamb/scale_ts1/genblk1[2].mult/added[2] ), 
        .C(n17691), .Y(n17667) );
  AOI21X1 U11420 ( .A(n17665), .B(n17664), .C(n18307), .Y(n18305) );
  INVX1 U11421 ( .A(n19753), .Y(n19752) );
  AND2X1 U11422 ( .A(n19752), .B(n18309), .Y(n18306) );
  INVX1 U11423 ( .A(n17666), .Y(n17770) );
  AOI21X1 U11424 ( .A(n16376), .B(n18306), .C(n17770), .Y(n17734) );
  INVX1 U11425 ( .A(n16985), .Y(n17703) );
  AOI21X1 U11426 ( .A(n17687), .B(n17667), .C(n17703), .Y(n17681) );
  OR2X1 U11427 ( .A(\lamb/scale_ds1/genblk1[2].mult/added[4] ), .B(
        \add_x_72/n1 ), .Y(n17718) );
  OR2X1 U11428 ( .A(n17718), .B(\lamb/scale_ds1/genblk1[2].mult/added[3] ), 
        .Y(n17674) );
  NAND2X1 U11429 ( .A(\lamb/scale_ds1/genblk1[2].mult/added[2] ), .B(n17674), 
        .Y(n17672) );
  INVX1 U11430 ( .A(n17672), .Y(n17669) );
  NAND2X1 U11431 ( .A(\lamb/scale_ds1/genblk1[2].mult/added[4] ), .B(
        \add_x_72/n1 ), .Y(n17670) );
  NAND3X1 U11432 ( .A(\lamb/scale_ds1/genblk1[2].mult/added[3] ), .B(n17670), 
        .C(n17718), .Y(n17719) );
  OR2X1 U11433 ( .A(\lamb/scale_ds1/genblk1[2].mult/added[1] ), .B(n17719), 
        .Y(n17710) );
  INVX1 U11434 ( .A(\lamb/scale_ds1/genblk1[2].mult/added[2] ), .Y(n17668) );
  NAND3X1 U11435 ( .A(\lamb/scale_ds1/genblk1[2].mult/added[4] ), .B(
        \add_x_72/n1 ), .C(\lamb/scale_ds1/genblk1[2].mult/added[3] ), .Y(
        n17677) );
  AOI22X1 U11436 ( .A(n17669), .B(n17710), .C(n17668), .D(n16586), .Y(n17684)
         );
  NAND2X1 U11437 ( .A(\lamb/scale_ds1/genblk1[2].mult/added[3] ), .B(n17718), 
        .Y(n17671) );
  INVX1 U11438 ( .A(\lamb/scale_ds1/genblk1[2].mult/added[3] ), .Y(n17717) );
  NAND2X1 U11439 ( .A(n17671), .B(n16999), .Y(n17673) );
  AOI22X1 U11440 ( .A(\lamb/scale_ds1/genblk1[2].mult/added[2] ), .B(
        \lamb/scale_ds1/genblk1[2].mult/added[1] ), .C(n17673), .D(n17672), 
        .Y(n17720) );
  INVX1 U11441 ( .A(n17720), .Y(n17678) );
  INVX1 U11442 ( .A(n17673), .Y(n17709) );
  INVX1 U11443 ( .A(n16586), .Y(n17676) );
  NAND2X1 U11444 ( .A(\lamb/scale_ds1/genblk1[2].mult/added[2] ), .B(
        \lamb/scale_ds1/genblk1[2].mult/added[1] ), .Y(n17675) );
  OAI21X1 U11445 ( .A(n17676), .B(n17675), .C(n17674), .Y(n17682) );
  AOI21X1 U11446 ( .A(\lamb/scale_ds1/genblk1[2].mult/added[1] ), .B(n17709), 
        .C(n17682), .Y(n17708) );
  OAI21X1 U11447 ( .A(n17678), .B(n16586), .C(n17708), .Y(n17679) );
  NAND2X1 U11448 ( .A(n18346), .B(n18344), .Y(n19721) );
  AOI21X1 U11449 ( .A(n19719), .B(n19721), .C(n18348), .Y(n19750) );
  AOI21X1 U11450 ( .A(n18346), .B(n16464), .C(n18344), .Y(n19749) );
  OAI21X1 U11451 ( .A(n17684), .B(n17679), .C(n17032), .Y(n17680) );
  HAX1 U11452 ( .A(n17681), .B(n17680), .YS(n19762) );
  OAI21X1 U11453 ( .A(n18334), .B(n17738), .C(n16419), .Y(n18029) );
  AOI22X1 U11454 ( .A(n18414), .B(n19762), .C(n18029), .D(n18412), .Y(n17740)
         );
  INVX1 U11455 ( .A(n17740), .Y(n17741) );
  INVX1 U11456 ( .A(\lamb/scale_ds1/genblk1[2].mult/added[1] ), .Y(n17707) );
  AOI21X1 U11457 ( .A(n17707), .B(n16999), .C(n17682), .Y(n17683) );
  OAI21X1 U11458 ( .A(n17684), .B(n17683), .C(n17032), .Y(n17693) );
  NAND2X1 U11459 ( .A(n17686), .B(n17685), .Y(n17732) );
  INVX1 U11460 ( .A(n17687), .Y(n17688) );
  AOI22X1 U11461 ( .A(n17689), .B(n17015), .C(n17732), .D(n17688), .Y(n17690)
         );
  OAI21X1 U11462 ( .A(n17691), .B(n17690), .C(n16985), .Y(n17692) );
  HAX1 U11463 ( .A(n17693), .B(n17692), .YS(n18245) );
  INVX1 U11464 ( .A(n18245), .Y(n18241) );
  NAND2X1 U11465 ( .A(n18336), .B(n17123), .Y(n17694) );
  OAI21X1 U11466 ( .A(n17695), .B(n18330), .C(n17694), .Y(n18202) );
  INVX1 U11467 ( .A(n18202), .Y(n18030) );
  AOI22X1 U11468 ( .A(n18414), .B(n18241), .C(n18030), .D(n18412), .Y(n17742)
         );
  AND2X1 U11469 ( .A(n17741), .B(n16590), .Y(n17749) );
  NAND3X1 U11470 ( .A(n17698), .B(n16941), .C(n16364), .Y(n17699) );
  OAI21X1 U11471 ( .A(\lamb/scale_ts1/genblk1[2].mult/added[2] ), .B(n16518), 
        .C(n17699), .Y(n17705) );
  NOR2X1 U11472 ( .A(n16458), .B(n17015), .Y(n17727) );
  NAND2X1 U11473 ( .A(n17727), .B(\lamb/scale_ts1/genblk1[2].mult/added[1] ), 
        .Y(n17704) );
  AOI21X1 U11474 ( .A(n17705), .B(n17704), .C(n17703), .Y(n17714) );
  NAND3X1 U11475 ( .A(\lamb/scale_ds1/genblk1[2].mult/added[2] ), .B(
        \lamb/scale_ds1/genblk1[2].mult/added[1] ), .C(n17706), .Y(n17724) );
  AOI22X1 U11476 ( .A(\lamb/scale_ds1/genblk1[2].mult/added[2] ), .B(n17709), 
        .C(n16961), .D(n17708), .Y(n17711) );
  NAND3X1 U11477 ( .A(n17724), .B(n17711), .C(n17710), .Y(n17712) );
  NAND2X1 U11478 ( .A(n17712), .B(n17032), .Y(n17713) );
  HAX1 U11479 ( .A(n17714), .B(n17713), .YS(n19765) );
  INVX1 U11480 ( .A(n19699), .Y(n18338) );
  NAND2X1 U11481 ( .A(n18338), .B(n17123), .Y(n17715) );
  OAI21X1 U11482 ( .A(n17716), .B(n16664), .C(n17715), .Y(n18205) );
  INVX1 U11483 ( .A(n18205), .Y(n19663) );
  AOI22X1 U11484 ( .A(n18414), .B(n19765), .C(n19663), .D(n18412), .Y(n17751)
         );
  INVX1 U11485 ( .A(n17094), .Y(n17745) );
  NAND2X1 U11486 ( .A(n17718), .B(n17717), .Y(n17721) );
  AOI22X1 U11487 ( .A(n16961), .B(n17721), .C(n17720), .D(n17719), .Y(n17725)
         );
  AOI21X1 U11488 ( .A(n17725), .B(n17724), .C(n17723), .Y(n17736) );
  INVX1 U11489 ( .A(n16320), .Y(n17728) );
  AOI22X1 U11490 ( .A(\lamb/scale_ts1/genblk1[2].mult/added[1] ), .B(n17728), 
        .C(\lamb/scale_ts1/genblk1[2].mult/added[2] ), .D(n17727), .Y(n17731)
         );
  INVX1 U11491 ( .A(n17729), .Y(n17730) );
  NAND3X1 U11492 ( .A(n17732), .B(n17731), .C(n17730), .Y(n17733) );
  NAND2X1 U11493 ( .A(n16985), .B(n17733), .Y(n17735) );
  HAX1 U11494 ( .A(n17736), .B(n17735), .YS(n19759) );
  NAND2X1 U11495 ( .A(n18337), .B(n17123), .Y(n17737) );
  OAI21X1 U11496 ( .A(n17739), .B(n16664), .C(n17737), .Y(n18206) );
  INVX1 U11497 ( .A(n18206), .Y(n18031) );
  AOI22X1 U11498 ( .A(n18414), .B(n19759), .C(n18031), .D(n18412), .Y(n17744)
         );
  OAI21X1 U11499 ( .A(n16334), .B(n17745), .C(n16599), .Y(
        \lamb/scale_ts3/genblk1[3].mult/logA[0] ) );
  INVX1 U11500 ( .A(n17744), .Y(n17750) );
  AND2X1 U11501 ( .A(n17750), .B(n17741), .Y(n19096) );
  AOI21X1 U11502 ( .A(n16590), .B(n16599), .C(n17094), .Y(n19095) );
  NOR3X1 U11503 ( .A(n19096), .B(n16372), .C(n17743), .Y(
        \lamb/scale_ts3/genblk1[3].mult/logA[1] ) );
  NAND2X1 U11504 ( .A(n17744), .B(n17094), .Y(n17754) );
  NOR2X1 U11505 ( .A(n17750), .B(n17018), .Y(n17746) );
  AOI22X1 U11506 ( .A(n17094), .B(n16599), .C(n17746), .D(n17745), .Y(n17748)
         );
  AOI21X1 U11507 ( .A(n17749), .B(n17754), .C(n17748), .Y(
        \lamb/scale_ts3/genblk1[3].mult/logA[2] ) );
  NAND2X1 U11508 ( .A(n17094), .B(n17750), .Y(n17752) );
  AOI22X1 U11509 ( .A(n17018), .B(n17754), .C(n16334), .D(n17752), .Y(
        \lamb/scale_ts3/genblk1[3].mult/logA[3] ) );
  INVX1 U11510 ( .A(\lamb/scale_ds1/genblk1[1].mult/added[3] ), .Y(n17759) );
  INVX1 U11511 ( .A(\lamb/scale_ds1/genblk1[1].mult/added[1] ), .Y(n17794) );
  INVX1 U11512 ( .A(n16503), .Y(n17789) );
  NAND2X1 U11513 ( .A(n17794), .B(n17789), .Y(n17758) );
  INVX1 U11514 ( .A(\lamb/scale_ds1/genblk1[1].mult/added[2] ), .Y(n17824) );
  NAND2X1 U11515 ( .A(n17789), .B(n16437), .Y(n17756) );
  OAI21X1 U11516 ( .A(n17776), .B(n17824), .C(n17756), .Y(n17757) );
  AOI22X1 U11517 ( .A(n16318), .B(n16354), .C(n17758), .D(n17757), .Y(n17760)
         );
  AOI21X1 U11518 ( .A(n17760), .B(n16906), .C(n16383), .Y(n17773) );
  OR2X1 U11519 ( .A(\lamb/scale_ts1/genblk1[1].mult/added[4] ), .B(
        \add_x_69/n1 ), .Y(n17798) );
  NOR2X1 U11520 ( .A(n17798), .B(\lamb/scale_ts1/genblk1[1].mult/added[3] ), 
        .Y(n17763) );
  INVX1 U11521 ( .A(n17798), .Y(n17761) );
  AOI21X1 U11522 ( .A(\add_x_69/n1 ), .B(
        \lamb/scale_ts1/genblk1[1].mult/added[4] ), .C(n17761), .Y(n17806) );
  INVX1 U11523 ( .A(\lamb/scale_ts1/genblk1[1].mult/added[1] ), .Y(n17816) );
  NAND3X1 U11524 ( .A(\lamb/scale_ts1/genblk1[1].mult/added[3] ), .B(n17010), 
        .C(n17816), .Y(n17809) );
  NAND3X1 U11525 ( .A(\lamb/scale_ts1/genblk1[1].mult/added[4] ), .B(
        \add_x_69/n1 ), .C(\lamb/scale_ts1/genblk1[1].mult/added[3] ), .Y(
        n17801) );
  INVX1 U11526 ( .A(\lamb/scale_ts1/genblk1[1].mult/added[2] ), .Y(n17800) );
  AOI22X1 U11527 ( .A(n17820), .B(n17809), .C(n16654), .D(n17800), .Y(n17783)
         );
  AND2X1 U11528 ( .A(\lamb/scale_ts1/genblk1[1].mult/added[4] ), .B(
        \add_x_69/n1 ), .Y(n17762) );
  NAND3X1 U11529 ( .A(n17762), .B(\lamb/scale_ts1/genblk1[1].mult/added[3] ), 
        .C(n17816), .Y(n17814) );
  NAND2X1 U11530 ( .A(\lamb/scale_ts1/genblk1[1].mult/added[1] ), .B(
        \lamb/scale_ts1/genblk1[1].mult/added[2] ), .Y(n17765) );
  INVX1 U11531 ( .A(n17765), .Y(n17764) );
  INVX1 U11532 ( .A(n17010), .Y(n17802) );
  NAND3X1 U11533 ( .A(n16945), .B(n16654), .C(n17802), .Y(n17815) );
  OR2X1 U11534 ( .A(\lamb/scale_ts1/genblk1[1].mult/added[3] ), .B(n17802), 
        .Y(n17819) );
  INVX1 U11535 ( .A(n17819), .Y(n17766) );
  AOI22X1 U11536 ( .A(\lamb/scale_ts1/genblk1[1].mult/added[1] ), .B(n16942), 
        .C(n17766), .D(n17765), .Y(n17785) );
  OR2X1 U11537 ( .A(n17815), .B(n17785), .Y(n17767) );
  NAND3X1 U11538 ( .A(n17814), .B(n16942), .C(n17767), .Y(n17771) );
  INVX1 U11539 ( .A(n19740), .Y(n18315) );
  AND2X1 U11540 ( .A(n18315), .B(n19743), .Y(n19748) );
  INVX1 U11541 ( .A(n18314), .Y(n18317) );
  AOI21X1 U11542 ( .A(n19743), .B(n18317), .C(n18315), .Y(n17769) );
  INVX1 U11543 ( .A(n17769), .Y(n19745) );
  AOI21X1 U11544 ( .A(n18317), .B(n19745), .C(n19746), .Y(n19744) );
  AOI21X1 U11545 ( .A(n19748), .B(n19744), .C(n17770), .Y(n17810) );
  OAI21X1 U11546 ( .A(n17783), .B(n17771), .C(n16319), .Y(n17772) );
  HAX1 U11547 ( .A(n17773), .B(n17772), .YS(n18260) );
  AOI22X1 U11548 ( .A(n18414), .B(n18260), .C(n16750), .D(n18412), .Y(n17835)
         );
  AOI22X1 U11549 ( .A(\lamb/scale_ds1/genblk1[1].mult/added[1] ), .B(n16318), 
        .C(n16631), .D(n16354), .Y(n17782) );
  AOI21X1 U11550 ( .A(n17789), .B(n17794), .C(
        \lamb/scale_ds1/genblk1[1].mult/added[2] ), .Y(n17779) );
  NAND3X1 U11551 ( .A(n16503), .B(n17794), .C(n17042), .Y(n17795) );
  NAND2X1 U11552 ( .A(n16906), .B(n17795), .Y(n17778) );
  MUX2X1 U11553 ( .B(n17779), .A(\lamb/scale_ds1/genblk1[1].mult/added[2] ), 
        .S(n17778), .Y(n17781) );
  AOI21X1 U11554 ( .A(n17782), .B(n17781), .C(n16383), .Y(n17787) );
  INVX1 U11555 ( .A(n17783), .Y(n17784) );
  INVX1 U11556 ( .A(n16319), .Y(n17821) );
  AOI21X1 U11557 ( .A(n17785), .B(n17784), .C(n17821), .Y(n17786) );
  HAX1 U11558 ( .A(n16879), .B(n17786), .YS(n18259) );
  INVX1 U11559 ( .A(n18259), .Y(n18254) );
  AOI22X1 U11560 ( .A(n18414), .B(n18254), .C(n16663), .D(n18412), .Y(n17842)
         );
  INVX1 U11561 ( .A(n16655), .Y(n17837) );
  AOI22X1 U11562 ( .A(n16758), .B(n17837), .C(n16655), .D(n16757), .Y(n17845)
         );
  NAND2X1 U11563 ( .A(n16437), .B(\lamb/scale_ds1/genblk1[1].mult/added[2] ), 
        .Y(n17791) );
  INVX1 U11564 ( .A(n17791), .Y(n17790) );
  AOI22X1 U11565 ( .A(\lamb/scale_ds1/genblk1[1].mult/added[1] ), .B(n16631), 
        .C(n17790), .D(n17789), .Y(n17796) );
  OAI21X1 U11566 ( .A(n16503), .B(\lamb/scale_ds1/genblk1[1].mult/added[2] ), 
        .C(n17791), .Y(n17793) );
  NAND3X1 U11567 ( .A(n17796), .B(n17831), .C(n17795), .Y(n17797) );
  NAND2X1 U11568 ( .A(\lamb/scale_ts1/genblk1[1].mult/added[3] ), .B(
        \lamb/scale_ts1/genblk1[1].mult/added[2] ), .Y(n17805) );
  INVX1 U11569 ( .A(n17805), .Y(n17799) );
  AOI22X1 U11570 ( .A(n17799), .B(n17798), .C(n17816), .D(n17017), .Y(n17804)
         );
  NAND2X1 U11571 ( .A(n16654), .B(n17800), .Y(n17803) );
  NAND3X1 U11572 ( .A(n17804), .B(n17803), .C(n17802), .Y(n17808) );
  NAND3X1 U11573 ( .A(n17010), .B(\lamb/scale_ts1/genblk1[1].mult/added[1] ), 
        .C(n17805), .Y(n17807) );
  NAND3X1 U11574 ( .A(n17809), .B(n17808), .C(n17807), .Y(n17811) );
  NAND2X1 U11575 ( .A(n17811), .B(n16319), .Y(n17812) );
  HAX1 U11576 ( .A(n16880), .B(n17812), .YS(n18262) );
  INVX1 U11577 ( .A(n18262), .Y(n18258) );
  AOI22X1 U11578 ( .A(n18414), .B(n18258), .C(n16761), .D(n18412), .Y(n17839)
         );
  INVX1 U11579 ( .A(n17815), .Y(n17817) );
  AOI22X1 U11580 ( .A(\lamb/scale_ts1/genblk1[1].mult/added[2] ), .B(n16822), 
        .C(n17817), .D(n17816), .Y(n17823) );
  NAND3X1 U11581 ( .A(\lamb/scale_ts1/genblk1[1].mult/added[1] ), .B(n17017), 
        .C(n17819), .Y(n17822) );
  AOI21X1 U11582 ( .A(n17823), .B(n17822), .C(n17821), .Y(n17833) );
  NAND2X1 U11583 ( .A(\lamb/scale_ds1/genblk1[1].mult/added[3] ), .B(n17824), 
        .Y(n17826) );
  AOI22X1 U11584 ( .A(n17776), .B(n17826), .C(
        \lamb/scale_ds1/genblk1[1].mult/added[2] ), .D(n16631), .Y(n17829) );
  OAI21X1 U11585 ( .A(\lamb/scale_ds1/genblk1[1].mult/added[1] ), .B(
        \lamb/scale_ds1/genblk1[1].mult/added[3] ), .C(n16629), .Y(n17828) );
  AOI22X1 U11586 ( .A(\lamb/scale_ds1/genblk1[1].mult/added[1] ), .B(
        \lamb/scale_ds1/genblk1[1].mult/added[2] ), .C(n17829), .D(n17828), 
        .Y(n17830) );
  OAI21X1 U11587 ( .A(n16895), .B(n17830), .C(n18369), .Y(n17832) );
  HAX1 U11588 ( .A(n17833), .B(n17832), .YS(n18261) );
  AOI22X1 U11589 ( .A(n18414), .B(n18261), .C(n16760), .D(n18412), .Y(n17843)
         );
  OAI21X1 U11590 ( .A(n16332), .B(n16742), .C(n16998), .Y(
        \lamb/scale_ts3/genblk1[2].mult/logA[0] ) );
  AOI21X1 U11591 ( .A(n16655), .B(n16998), .C(n16743), .Y(n18971) );
  NOR3X1 U11592 ( .A(n16758), .B(n16742), .C(n17837), .Y(n17834) );
  NOR3X1 U11593 ( .A(n16368), .B(n16373), .C(n17834), .Y(
        \lamb/scale_ts3/genblk1[2].mult/logA[1] ) );
  NOR2X1 U11594 ( .A(n17837), .B(n16758), .Y(n17841) );
  NAND2X1 U11595 ( .A(n16747), .B(n16743), .Y(n17846) );
  OAI21X1 U11596 ( .A(n16743), .B(n17837), .C(n17836), .Y(n17838) );
  OAI21X1 U11597 ( .A(n16743), .B(n16747), .C(n17838), .Y(n17840) );
  AOI21X1 U11598 ( .A(n17841), .B(n17846), .C(n17840), .Y(
        \lamb/scale_ts3/genblk1[2].mult/logA[2] ) );
  OR2X1 U11599 ( .A(n16742), .B(n16747), .Y(n17844) );
  AOI22X1 U11600 ( .A(n16823), .B(n17846), .C(n16332), .D(n17844), .Y(
        \lamb/scale_ts3/genblk1[2].mult/logA[3] ) );
  NAND3X1 U11601 ( .A(\add_x_59/n1 ), .B(
        \lamb/scale_ds2/genblk1[2].mult/added[4] ), .C(
        \lamb/scale_ds2/genblk1[2].mult/added[3] ), .Y(n17900) );
  INVX1 U11602 ( .A(n16646), .Y(n17849) );
  NAND2X1 U11603 ( .A(\lamb/scale_ds2/genblk1[2].mult/added[1] ), .B(
        \lamb/scale_ds2/genblk1[2].mult/added[2] ), .Y(n17848) );
  OR2X1 U11604 ( .A(\add_x_59/n1 ), .B(
        \lamb/scale_ds2/genblk1[2].mult/added[4] ), .Y(n17864) );
  OR2X1 U11605 ( .A(n17864), .B(\lamb/scale_ds2/genblk1[2].mult/added[3] ), 
        .Y(n17852) );
  OAI21X1 U11606 ( .A(n17849), .B(n17848), .C(n17852), .Y(n17865) );
  AOI21X1 U11607 ( .A(\lamb/scale_ds2/genblk1[2].mult/added[4] ), .B(
        \add_x_59/n1 ), .C(\lamb/scale_ds2/genblk1[2].mult/added[3] ), .Y(
        n17880) );
  NAND2X1 U11608 ( .A(\lamb/scale_ds2/genblk1[2].mult/added[3] ), .B(n17864), 
        .Y(n17883) );
  INVX1 U11609 ( .A(n17883), .Y(n17851) );
  NOR2X1 U11610 ( .A(n16530), .B(n17851), .Y(n17879) );
  INVX1 U11611 ( .A(n17879), .Y(n17902) );
  INVX1 U11612 ( .A(\lamb/scale_ds2/genblk1[2].mult/added[1] ), .Y(n17901) );
  OAI21X1 U11613 ( .A(n17902), .B(n17901), .C(n16646), .Y(n17854) );
  NAND2X1 U11614 ( .A(\add_x_59/n1 ), .B(
        \lamb/scale_ds2/genblk1[2].mult/added[4] ), .Y(n17850) );
  NAND3X1 U11615 ( .A(n17851), .B(n17850), .C(n17901), .Y(n17881) );
  NAND3X1 U11616 ( .A(n17852), .B(n16966), .C(
        \lamb/scale_ds2/genblk1[2].mult/added[2] ), .Y(n17853) );
  OAI21X1 U11617 ( .A(\lamb/scale_ds2/genblk1[2].mult/added[2] ), .B(n17854), 
        .C(n17853), .Y(n17868) );
  OAI21X1 U11618 ( .A(\lamb/scale_ds2/genblk1[2].mult/added[1] ), .B(n16646), 
        .C(n17868), .Y(n17856) );
  INVX1 U11619 ( .A(n18260), .Y(n18250) );
  NAND3X1 U11620 ( .A(n18254), .B(n18258), .C(n18261), .Y(n17855) );
  OR2X1 U11621 ( .A(n18250), .B(n17855), .Y(n17884) );
  OAI21X1 U11622 ( .A(n17865), .B(n17856), .C(n17884), .Y(n17863) );
  NAND2X1 U11623 ( .A(\lamb/scale_ts2/genblk1[2].mult/added[4] ), .B(
        \add_x_55/n1 ), .Y(n17914) );
  INVX1 U11624 ( .A(n17914), .Y(n17891) );
  OR2X1 U11625 ( .A(n17891), .B(n16749), .Y(n17894) );
  NAND2X1 U11626 ( .A(\lamb/scale_ts2/genblk1[2].mult/added[3] ), .B(
        \lamb/scale_ts2/genblk1[2].mult/added[2] ), .Y(n17888) );
  INVX1 U11627 ( .A(n17888), .Y(n17889) );
  NAND3X1 U11628 ( .A(\lamb/scale_ts2/genblk1[2].mult/added[4] ), .B(
        \add_x_55/n1 ), .C(\lamb/scale_ts2/genblk1[2].mult/added[3] ), .Y(
        n17869) );
  INVX1 U11629 ( .A(\lamb/scale_ts2/genblk1[2].mult/added[3] ), .Y(n17873) );
  NAND2X1 U11630 ( .A(n16749), .B(n17873), .Y(n17857) );
  AOI22X1 U11631 ( .A(n16362), .B(n17889), .C(n16920), .D(n16369), .Y(n17861)
         );
  INVX1 U11632 ( .A(n17894), .Y(n17917) );
  INVX1 U11633 ( .A(\lamb/scale_ts2/genblk1[2].mult/added[2] ), .Y(n17870) );
  NAND2X1 U11634 ( .A(n17917), .B(n17870), .Y(n17858) );
  NAND3X1 U11635 ( .A(\lamb/scale_ts2/genblk1[2].mult/added[1] ), .B(n16589), 
        .C(n17858), .Y(n17860) );
  OAI21X1 U11636 ( .A(n16650), .B(n16663), .C(n16761), .Y(n18213) );
  NAND2X1 U11637 ( .A(n16760), .B(n18221), .Y(n17859) );
  OAI21X1 U11638 ( .A(n18213), .B(n17859), .C(n16619), .Y(n17919) );
  AOI21X1 U11639 ( .A(n17861), .B(n17860), .C(n17919), .Y(n17862) );
  HAX1 U11640 ( .A(n17863), .B(n17862), .YS(n17933) );
  INVX1 U11641 ( .A(n17933), .Y(n17925) );
  AOI21X1 U11642 ( .A(n17063), .B(n17901), .C(n17865), .Y(n17866) );
  INVX1 U11643 ( .A(n17866), .Y(n17867) );
  INVX1 U11644 ( .A(n17884), .Y(n17906) );
  AOI21X1 U11645 ( .A(n17868), .B(n17867), .C(n17906), .Y(n17878) );
  AOI22X1 U11646 ( .A(\lamb/scale_ts2/genblk1[2].mult/added[2] ), .B(n16589), 
        .C(n16749), .D(n17873), .Y(n17872) );
  AOI22X1 U11647 ( .A(n17872), .B(\lamb/scale_ts2/genblk1[2].mult/added[1] ), 
        .C(n16362), .D(n17050), .Y(n17876) );
  NAND2X1 U11648 ( .A(n17050), .B(n16321), .Y(n17874) );
  NAND2X1 U11649 ( .A(n16920), .B(n17874), .Y(n17887) );
  AOI21X1 U11650 ( .A(n17876), .B(n17887), .C(n17919), .Y(n17877) );
  HAX1 U11651 ( .A(n16877), .B(n17877), .YS(n17932) );
  INVX1 U11652 ( .A(n17932), .Y(n17927) );
  AOI22X1 U11653 ( .A(n17925), .B(n17927), .C(n17932), .D(n17933), .Y(n17937)
         );
  AOI22X1 U11654 ( .A(n17903), .B(\lamb/scale_ds2/genblk1[2].mult/added[1] ), 
        .C(\lamb/scale_ds2/genblk1[2].mult/added[2] ), .D(n17879), .Y(n17882)
         );
  NAND3X1 U11655 ( .A(n16530), .B(\lamb/scale_ds2/genblk1[2].mult/added[1] ), 
        .C(\lamb/scale_ds2/genblk1[2].mult/added[2] ), .Y(n17907) );
  NAND3X1 U11656 ( .A(n17882), .B(n17907), .C(n16966), .Y(n17886) );
  NOR3X1 U11657 ( .A(\lamb/scale_ds2/genblk1[2].mult/added[2] ), .B(n17901), 
        .C(n17883), .Y(n17885) );
  OAI21X1 U11658 ( .A(n17886), .B(n17885), .C(n17884), .Y(n17899) );
  INVX1 U11659 ( .A(\lamb/scale_ts2/genblk1[2].mult/added[1] ), .Y(n17910) );
  OR2X1 U11660 ( .A(n17887), .B(n17910), .Y(n17920) );
  INVX1 U11661 ( .A(n17920), .Y(n17897) );
  AOI22X1 U11662 ( .A(\lamb/scale_ts2/genblk1[2].mult/added[1] ), .B(n17888), 
        .C(\lamb/scale_ts2/genblk1[2].mult/added[3] ), .D(n17910), .Y(n17893)
         );
  INVX1 U11663 ( .A(n16321), .Y(n17890) );
  AOI22X1 U11664 ( .A(n17891), .B(n17890), .C(n16749), .D(n17889), .Y(n17892)
         );
  OAI21X1 U11665 ( .A(n17894), .B(n17893), .C(n16794), .Y(n17896) );
  INVX1 U11666 ( .A(n17919), .Y(n17895) );
  OAI21X1 U11667 ( .A(n17897), .B(n17896), .C(n17895), .Y(n17898) );
  HAX1 U11668 ( .A(n17899), .B(n17898), .YS(n17929) );
  INVX1 U11669 ( .A(n17929), .Y(n17935) );
  AOI21X1 U11670 ( .A(n17063), .B(n16646), .C(
        \lamb/scale_ds2/genblk1[2].mult/added[1] ), .Y(n17905) );
  AOI22X1 U11671 ( .A(\lamb/scale_ds2/genblk1[2].mult/added[1] ), .B(
        \lamb/scale_ds2/genblk1[2].mult/added[2] ), .C(n17902), .D(n17901), 
        .Y(n17904) );
  AOI22X1 U11672 ( .A(n17905), .B(\lamb/scale_ds2/genblk1[2].mult/added[2] ), 
        .C(n17904), .D(n17063), .Y(n17908) );
  AOI21X1 U11673 ( .A(n17908), .B(n17907), .C(n17906), .Y(n17923) );
  OAI21X1 U11674 ( .A(n17050), .B(n17910), .C(n16321), .Y(n17918) );
  OAI21X1 U11675 ( .A(\lamb/scale_ts2/genblk1[2].mult/added[3] ), .B(
        \lamb/scale_ts2/genblk1[2].mult/added[1] ), .C(n16749), .Y(n17913) );
  OAI21X1 U11676 ( .A(n17911), .B(n17914), .C(n17913), .Y(n17915) );
  AOI22X1 U11677 ( .A(n17918), .B(n17917), .C(n16369), .D(n17915), .Y(n17921)
         );
  AOI21X1 U11678 ( .A(n17921), .B(n17920), .C(n17919), .Y(n17922) );
  HAX1 U11679 ( .A(n17923), .B(n17922), .YS(n17934) );
  OAI21X1 U11680 ( .A(n17937), .B(n17935), .C(n16997), .Y(
        \lamb/scale_ds3/genblk1[3].mult/logA[0] ) );
  NOR2X1 U11681 ( .A(n17934), .B(n17925), .Y(n19106) );
  AOI21X1 U11682 ( .A(n17932), .B(n16997), .C(n17929), .Y(n19105) );
  NOR3X1 U11683 ( .A(n17925), .B(n17927), .C(n17935), .Y(n17924) );
  NOR3X1 U11684 ( .A(n19106), .B(n19105), .C(n17924), .Y(
        \lamb/scale_ds3/genblk1[3].mult/logA[1] ) );
  NOR2X1 U11685 ( .A(n17927), .B(n17925), .Y(n17931) );
  NAND2X1 U11686 ( .A(n17934), .B(n17929), .Y(n17938) );
  OAI21X1 U11687 ( .A(n17929), .B(n17927), .C(n17926), .Y(n17928) );
  OAI21X1 U11688 ( .A(n17929), .B(n17934), .C(n17928), .Y(n17930) );
  AOI21X1 U11689 ( .A(n17931), .B(n17938), .C(n17930), .Y(
        \lamb/scale_ds3/genblk1[3].mult/logA[2] ) );
  NOR2X1 U11690 ( .A(n17933), .B(n17932), .Y(n17939) );
  OR2X1 U11691 ( .A(n17935), .B(n17934), .Y(n17936) );
  NAND3X1 U11692 ( .A(\lamb/scale_ts2/genblk1[1].mult/added[3] ), .B(
        \lamb/scale_ts2/genblk1[1].mult/added[4] ), .C(\add_x_56/n1 ), .Y(
        n17940) );
  NAND2X1 U11693 ( .A(\lamb/scale_ts2/genblk1[1].mult/added[2] ), .B(n17940), 
        .Y(n17980) );
  NAND2X1 U11694 ( .A(\lamb/scale_ts2/genblk1[1].mult/added[4] ), .B(
        \add_x_56/n1 ), .Y(n17941) );
  OR2X1 U11695 ( .A(\lamb/scale_ts2/genblk1[1].mult/added[4] ), .B(
        \add_x_56/n1 ), .Y(n17942) );
  INVX1 U11696 ( .A(n17941), .Y(n17944) );
  OR2X1 U11697 ( .A(\lamb/scale_ts2/genblk1[1].mult/added[3] ), .B(n17944), 
        .Y(n18003) );
  NOR2X1 U11698 ( .A(n17942), .B(\lamb/scale_ts2/genblk1[1].mult/added[3] ), 
        .Y(n17979) );
  INVX1 U11699 ( .A(n17979), .Y(n18004) );
  AND2X1 U11700 ( .A(\lamb/scale_ts2/genblk1[1].mult/added[2] ), .B(
        \lamb/scale_ts2/genblk1[1].mult/added[3] ), .Y(n17943) );
  INVX1 U11701 ( .A(\lamb/scale_ts2/genblk1[1].mult/added[1] ), .Y(n18001) );
  NAND3X1 U11702 ( .A(n17943), .B(n17942), .C(n18001), .Y(n17945) );
  INVX1 U11703 ( .A(\lamb/scale_ts2/genblk1[1].mult/added[2] ), .Y(n17977) );
  NAND3X1 U11704 ( .A(\lamb/scale_ts2/genblk1[1].mult/added[3] ), .B(n17944), 
        .C(n17977), .Y(n17982) );
  NAND3X1 U11705 ( .A(n18004), .B(n17945), .C(n16967), .Y(n17946) );
  AOI21X1 U11706 ( .A(\lamb/scale_ts2/genblk1[1].mult/added[1] ), .B(n16816), 
        .C(n17946), .Y(n17959) );
  AOI21X1 U11707 ( .A(n17950), .B(n17949), .C(n17948), .Y(n18008) );
  INVX1 U11708 ( .A(n16649), .Y(n17958) );
  INVX1 U11709 ( .A(\lamb/scale_ds2/genblk1[1].mult/added[3] ), .Y(n17966) );
  OAI21X1 U11710 ( .A(\lamb/scale_ds2/genblk1[1].mult/added[3] ), .B(
        \lamb/scale_ds2/genblk1[1].mult/added[1] ), .C(n17045), .Y(n17951) );
  NOR2X1 U11711 ( .A(n16324), .B(n17951), .Y(n17972) );
  NAND2X1 U11712 ( .A(n17972), .B(\lamb/scale_ds2/genblk1[1].mult/added[2] ), 
        .Y(n17990) );
  AOI21X1 U11713 ( .A(n17985), .B(n17990), .C(
        \lamb/scale_ds2/genblk1[1].mult/added[1] ), .Y(n17956) );
  INVX1 U11714 ( .A(\lamb/scale_ds2/genblk1[1].mult/added[2] ), .Y(n17984) );
  INVX1 U11715 ( .A(n17985), .Y(n17964) );
  INVX1 U11716 ( .A(n16324), .Y(n17967) );
  OAI21X1 U11717 ( .A(n17967), .B(n17966), .C(n17045), .Y(n18000) );
  OAI21X1 U11718 ( .A(n18000), .B(\lamb/scale_ds2/genblk1[1].mult/added[2] ), 
        .C(\lamb/scale_ds2/genblk1[1].mult/added[1] ), .Y(n17953) );
  OAI21X1 U11719 ( .A(n17964), .B(n17953), .C(n17009), .Y(n17954) );
  AOI21X1 U11720 ( .A(n17984), .B(n17964), .C(n17954), .Y(n17971) );
  INVX1 U11721 ( .A(n17971), .Y(n17955) );
  OAI21X1 U11722 ( .A(n17956), .B(n17955), .C(n18278), .Y(n17957) );
  OAI21X1 U11723 ( .A(n17959), .B(n17958), .C(n17957), .Y(n18018) );
  INVX1 U11724 ( .A(n18018), .Y(n18022) );
  AND2X1 U11725 ( .A(n18001), .B(n17960), .Y(n17978) );
  AOI22X1 U11726 ( .A(\lamb/scale_ts2/genblk1[1].mult/added[2] ), .B(
        \lamb/scale_ts2/genblk1[1].mult/added[3] ), .C(n17961), .D(n17977), 
        .Y(n17962) );
  AOI22X1 U11727 ( .A(\lamb/scale_ts2/genblk1[1].mult/added[3] ), .B(n17978), 
        .C(\lamb/scale_ts2/genblk1[1].mult/added[1] ), .D(n17962), .Y(n17963)
         );
  OAI21X1 U11728 ( .A(n17977), .B(n16600), .C(n17963), .Y(n17976) );
  INVX1 U11729 ( .A(n18000), .Y(n17974) );
  AOI22X1 U11730 ( .A(\lamb/scale_ds2/genblk1[1].mult/added[2] ), .B(
        \lamb/scale_ds2/genblk1[1].mult/added[1] ), .C(n17964), .D(n17984), 
        .Y(n17999) );
  INVX1 U11731 ( .A(n17999), .Y(n17970) );
  NAND3X1 U11732 ( .A(n17045), .B(n17967), .C(n17966), .Y(n17991) );
  NAND2X1 U11733 ( .A(\lamb/scale_ds2/genblk1[1].mult/added[2] ), .B(n17009), 
        .Y(n17986) );
  NAND2X1 U11734 ( .A(n17967), .B(n17966), .Y(n17968) );
  NAND3X1 U11735 ( .A(\lamb/scale_ds2/genblk1[1].mult/added[1] ), .B(n17986), 
        .C(n17968), .Y(n17969) );
  OAI21X1 U11736 ( .A(n17991), .B(n17984), .C(n17969), .Y(n17998) );
  AOI22X1 U11737 ( .A(n17972), .B(n17971), .C(n17970), .D(n17998), .Y(n17973)
         );
  OAI21X1 U11738 ( .A(n17974), .B(n16374), .C(n17973), .Y(n17975) );
  AOI22X1 U11739 ( .A(n16649), .B(n17976), .C(n18278), .D(n17975), .Y(n19708)
         );
  AOI22X1 U11740 ( .A(\lamb/scale_ts2/genblk1[1].mult/added[2] ), .B(n17979), 
        .C(n17978), .D(n16337), .Y(n17983) );
  NAND3X1 U11741 ( .A(\lamb/scale_ts2/genblk1[1].mult/added[1] ), .B(n18004), 
        .C(n17980), .Y(n17981) );
  NAND3X1 U11742 ( .A(n17983), .B(n16967), .C(n17981), .Y(n17997) );
  NAND2X1 U11743 ( .A(n16796), .B(n17986), .Y(n17995) );
  NAND3X1 U11744 ( .A(\lamb/scale_ds2/genblk1[1].mult/added[1] ), .B(n17009), 
        .C(n16374), .Y(n17994) );
  AOI21X1 U11745 ( .A(n17991), .B(n17990), .C(
        \lamb/scale_ds2/genblk1[1].mult/added[1] ), .Y(n17992) );
  INVX1 U11746 ( .A(n17992), .Y(n17993) );
  NAND3X1 U11747 ( .A(n17995), .B(n17994), .C(n17993), .Y(n17996) );
  AOI22X1 U11748 ( .A(n16649), .B(n17997), .C(n18278), .D(n17996), .Y(n18019)
         );
  AOI21X1 U11749 ( .A(n18000), .B(n17999), .C(n17998), .Y(n18012) );
  AOI21X1 U11750 ( .A(n18004), .B(n16337), .C(n18001), .Y(n18010) );
  OAI21X1 U11751 ( .A(n17960), .B(\lamb/scale_ts2/genblk1[1].mult/added[1] ), 
        .C(n18003), .Y(n18005) );
  NAND3X1 U11752 ( .A(n18005), .B(n18004), .C(
        \lamb/scale_ts2/genblk1[1].mult/added[2] ), .Y(n18006) );
  OAI21X1 U11753 ( .A(\lamb/scale_ts2/genblk1[1].mult/added[2] ), .B(n16600), 
        .C(n18006), .Y(n18009) );
  OAI21X1 U11754 ( .A(n16818), .B(n18009), .C(n16649), .Y(n18011) );
  OAI21X1 U11755 ( .A(n18012), .B(n16479), .C(n18011), .Y(n18020) );
  OAI21X1 U11756 ( .A(n17080), .B(n16632), .C(n18020), .Y(n18013) );
  INVX1 U11757 ( .A(n16632), .Y(n18021) );
  INVX1 U11758 ( .A(n17080), .Y(n18014) );
  AOI21X1 U11759 ( .A(n16598), .B(n18021), .C(n18014), .Y(n18985) );
  AOI21X1 U11760 ( .A(n18022), .B(n18013), .C(n18985), .Y(
        \lamb/scale_ds3/genblk1[2].mult/logA[1] ) );
  INVX1 U11761 ( .A(n18020), .Y(n18017) );
  AOI21X1 U11762 ( .A(n18014), .B(n18020), .C(n16632), .Y(n18015) );
  MUX2X1 U11763 ( .B(n16598), .A(n18018), .S(n18015), .Y(n18016) );
  AOI21X1 U11764 ( .A(n17080), .B(n18017), .C(n18016), .Y(
        \lamb/scale_ds3/genblk1[2].mult/logA[2] ) );
  NOR2X1 U11765 ( .A(n18020), .B(n19705), .Y(n18984) );
  AOI21X1 U11766 ( .A(n19705), .B(n18020), .C(n18984), .Y(n18023) );
  NAND2X1 U11767 ( .A(n18022), .B(n18021), .Y(n19704) );
  OAI21X1 U11768 ( .A(n17080), .B(n18023), .C(n19704), .Y(
        \lamb/scale_ds3/genblk1[2].mult/logA[3] ) );
  NOR3X1 U11769 ( .A(\lamb/scale_ts2/genblk1[3].mult/added[3] ), .B(
        \lamb/scale_ts2/genblk1[3].mult/added[4] ), .C(\add_x_54/n1 ), .Y(
        n18026) );
  NOR2X1 U11770 ( .A(\lamb/scale_ts2/genblk1[3].mult/added[4] ), .B(
        \add_x_54/n1 ), .Y(n18068) );
  INVX1 U11771 ( .A(n18068), .Y(n18082) );
  AOI21X1 U11772 ( .A(\lamb/scale_ts2/genblk1[3].mult/added[4] ), .B(
        \add_x_54/n1 ), .C(n16572), .Y(n18047) );
  INVX1 U11773 ( .A(\lamb/scale_ts2/genblk1[3].mult/added[1] ), .Y(n18086) );
  NAND2X1 U11774 ( .A(n18047), .B(n18086), .Y(n18073) );
  INVX1 U11775 ( .A(n18073), .Y(n18024) );
  OAI21X1 U11776 ( .A(n18026), .B(n18024), .C(
        \lamb/scale_ts2/genblk1[3].mult/added[2] ), .Y(n18033) );
  AND2X1 U11777 ( .A(\lamb/scale_ts2/genblk1[3].mult/added[4] ), .B(
        \add_x_54/n1 ), .Y(n18025) );
  OR2X1 U11778 ( .A(\lamb/scale_ts2/genblk1[3].mult/added[3] ), .B(n18025), 
        .Y(n18070) );
  OAI21X1 U11779 ( .A(\lamb/scale_ts2/genblk1[3].mult/added[2] ), .B(n17048), 
        .C(n18070), .Y(n18027) );
  INVX1 U11780 ( .A(\lamb/scale_ts2/genblk1[3].mult/added[2] ), .Y(n18084) );
  NOR2X1 U11781 ( .A(n18086), .B(n18084), .Y(n18049) );
  OAI21X1 U11782 ( .A(n18026), .B(n18049), .C(n17048), .Y(n18046) );
  OAI21X1 U11783 ( .A(\lamb/scale_ts2/genblk1[3].mult/added[1] ), .B(n18027), 
        .C(n18046), .Y(n18032) );
  NAND2X1 U11784 ( .A(n18205), .B(n18202), .Y(n18028) );
  INVX1 U11785 ( .A(n18029), .Y(n18198) );
  AOI21X1 U11786 ( .A(n18206), .B(n18028), .C(n18198), .Y(n18199) );
  NAND2X1 U11787 ( .A(n18198), .B(n18030), .Y(n18208) );
  NAND2X1 U11788 ( .A(n16888), .B(n18208), .Y(n19660) );
  AOI21X1 U11789 ( .A(n18031), .B(n18205), .C(n19660), .Y(n18209) );
  AOI21X1 U11790 ( .A(n18199), .B(n18209), .C(n17948), .Y(n18075) );
  INVX1 U11791 ( .A(n16984), .Y(n18087) );
  AOI21X1 U11792 ( .A(n18033), .B(n18032), .C(n18087), .Y(n18045) );
  INVX1 U11793 ( .A(\lamb/scale_ds2/genblk1[3].mult/added[1] ), .Y(n18053) );
  AND2X1 U11794 ( .A(\lamb/scale_ds2/genblk1[3].mult/added[2] ), .B(n18053), 
        .Y(n18036) );
  AND2X1 U11795 ( .A(\lamb/scale_ds2/genblk1[3].mult/added[4] ), .B(
        \add_x_58/n1 ), .Y(n18034) );
  INVX1 U11796 ( .A(\lamb/scale_ds2/genblk1[3].mult/added[3] ), .Y(n18056) );
  NOR3X1 U11797 ( .A(n18034), .B(n17041), .C(n18056), .Y(n18064) );
  NAND3X1 U11798 ( .A(\lamb/scale_ds2/genblk1[3].mult/added[4] ), .B(
        \add_x_58/n1 ), .C(\lamb/scale_ds2/genblk1[3].mult/added[3] ), .Y(
        n18039) );
  NAND2X1 U11799 ( .A(\lamb/scale_ds2/genblk1[3].mult/added[2] ), .B(n17041), 
        .Y(n18035) );
  AOI22X1 U11800 ( .A(\lamb/scale_ds2/genblk1[3].mult/added[2] ), .B(
        \lamb/scale_ds2/genblk1[3].mult/added[3] ), .C(n18039), .D(n18035), 
        .Y(n18063) );
  AOI21X1 U11801 ( .A(n18036), .B(n18064), .C(n18063), .Y(n18037) );
  INVX1 U11802 ( .A(n18037), .Y(n18060) );
  NAND2X1 U11803 ( .A(n18056), .B(n18038), .Y(n18094) );
  AOI21X1 U11804 ( .A(\lamb/scale_ds2/genblk1[3].mult/added[4] ), .B(
        \add_x_58/n1 ), .C(n18094), .Y(n18092) );
  INVX1 U11805 ( .A(n16573), .Y(n18041) );
  NAND2X1 U11806 ( .A(n17041), .B(n18056), .Y(n18040) );
  INVX1 U11807 ( .A(n18039), .Y(n18054) );
  AOI21X1 U11808 ( .A(n16630), .B(n18040), .C(n18054), .Y(n18052) );
  AOI21X1 U11809 ( .A(n18053), .B(n18041), .C(n18052), .Y(n18043) );
  NAND2X1 U11810 ( .A(n19759), .B(n19762), .Y(n18246) );
  NAND2X1 U11811 ( .A(n18241), .B(n19765), .Y(n18042) );
  OR2X1 U11812 ( .A(n18246), .B(n18042), .Y(n18098) );
  OAI21X1 U11813 ( .A(n18060), .B(n16830), .C(n18098), .Y(n18044) );
  HAX1 U11814 ( .A(n18045), .B(n18044), .YS(n18407) );
  INVX1 U11815 ( .A(n18407), .Y(n19776) );
  INVX1 U11816 ( .A(n18046), .Y(n18051) );
  AOI22X1 U11817 ( .A(\lamb/scale_ts2/genblk1[3].mult/added[1] ), .B(n18081), 
        .C(n18047), .D(\lamb/scale_ts2/genblk1[3].mult/added[2] ), .Y(n18048)
         );
  OAI21X1 U11818 ( .A(n18049), .B(n17048), .C(n18048), .Y(n18050) );
  OAI21X1 U11819 ( .A(n18051), .B(n18050), .C(n16984), .Y(n18062) );
  INVX1 U11820 ( .A(n18052), .Y(n18058) );
  NAND3X1 U11821 ( .A(n18054), .B(\lamb/scale_ds2/genblk1[3].mult/added[2] ), 
        .C(n18053), .Y(n18097) );
  NAND3X1 U11822 ( .A(\add_x_58/n1 ), .B(
        \lamb/scale_ds2/genblk1[3].mult/added[4] ), .C(n18056), .Y(n18055) );
  OAI21X1 U11823 ( .A(n18038), .B(n18056), .C(n18055), .Y(n18090) );
  NAND2X1 U11824 ( .A(\lamb/scale_ds2/genblk1[3].mult/added[1] ), .B(n18090), 
        .Y(n18057) );
  OAI21X1 U11825 ( .A(n18060), .B(n18059), .C(n18098), .Y(n18061) );
  HAX1 U11826 ( .A(n18062), .B(n18061), .YS(n18104) );
  INVX1 U11827 ( .A(n18104), .Y(n19778) );
  AOI22X1 U11828 ( .A(n19776), .B(n19778), .C(n18104), .D(n18407), .Y(n18106)
         );
  OAI21X1 U11829 ( .A(n16573), .B(n18063), .C(
        \lamb/scale_ds2/genblk1[3].mult/added[1] ), .Y(n18067) );
  AOI22X1 U11830 ( .A(\lamb/scale_ds2/genblk1[3].mult/added[2] ), .B(n18090), 
        .C(n18064), .D(n16630), .Y(n18066) );
  INVX1 U11831 ( .A(n18098), .Y(n18065) );
  AOI21X1 U11832 ( .A(n18067), .B(n18066), .C(n18065), .Y(n18077) );
  NOR2X1 U11833 ( .A(n18070), .B(n18068), .Y(n18079) );
  AOI22X1 U11834 ( .A(\lamb/scale_ts2/genblk1[3].mult/added[1] ), .B(n18079), 
        .C(\lamb/scale_ts2/genblk1[3].mult/added[2] ), .D(n18081), .Y(n18072)
         );
  MUX2X1 U11835 ( .B(n18070), .A(n16572), .S(n18084), .Y(n18071) );
  NAND3X1 U11836 ( .A(n18073), .B(n18072), .C(n16963), .Y(n18074) );
  NAND2X1 U11837 ( .A(n16984), .B(n18074), .Y(n18076) );
  HAX1 U11838 ( .A(n18077), .B(n18076), .YS(n19775) );
  OAI21X1 U11839 ( .A(n18079), .B(n18078), .C(
        \lamb/scale_ts2/genblk1[3].mult/added[2] ), .Y(n18080) );
  NAND2X1 U11840 ( .A(n16986), .B(n18080), .Y(n18085) );
  OAI21X1 U11841 ( .A(n18086), .B(n18082), .C(n16986), .Y(n18083) );
  AOI22X1 U11842 ( .A(n18086), .B(n18085), .C(n18084), .D(n18083), .Y(n18088)
         );
  AOI21X1 U11843 ( .A(n16963), .B(n18088), .C(n18087), .Y(n18101) );
  AOI22X1 U11844 ( .A(\lamb/scale_ds2/genblk1[3].mult/added[2] ), .B(n16573), 
        .C(n16630), .D(n18090), .Y(n18096) );
  NAND2X1 U11845 ( .A(\lamb/scale_ds2/genblk1[3].mult/added[3] ), .B(
        \lamb/scale_ds2/genblk1[3].mult/added[2] ), .Y(n18093) );
  NAND3X1 U11846 ( .A(\lamb/scale_ds2/genblk1[3].mult/added[1] ), .B(n18094), 
        .C(n18093), .Y(n18095) );
  NAND3X1 U11847 ( .A(n18097), .B(n18096), .C(n18095), .Y(n18099) );
  XNOR2X1 U11848 ( .A(n18101), .B(n16881), .Y(n18405) );
  OAI21X1 U11849 ( .A(n16333), .B(n19775), .C(n16407), .Y(
        \lamb/scale_bs3/genblk1[0].mult/logB[0] ) );
  OAI21X1 U11850 ( .A(n18407), .B(n19775), .C(n18405), .Y(n18103) );
  NAND2X1 U11851 ( .A(n19776), .B(n16407), .Y(n18102) );
  AOI22X1 U11852 ( .A(n19778), .B(n18103), .C(n19775), .D(n18102), .Y(
        \lamb/scale_bs3/genblk1[0].mult/logB[1] ) );
  AND2X1 U11853 ( .A(n18407), .B(n18104), .Y(n18107) );
  INVX1 U11854 ( .A(n19775), .Y(n18406) );
  OR2X1 U11855 ( .A(n19775), .B(n18405), .Y(n18105) );
  AOI22X1 U11856 ( .A(n18107), .B(n16325), .C(n16333), .D(n18105), .Y(
        \lamb/scale_bs3/genblk1[0].mult/logB[3] ) );
  INVX1 U11857 ( .A(\lamb/scale_ls2/genblk1[2].mult/added[1] ), .Y(n18109) );
  AND2X1 U11858 ( .A(\lamb/scale_ls2/genblk1[2].mult/added[3] ), .B(n18114), 
        .Y(n19733) );
  NAND2X1 U11859 ( .A(\lamb/scale_ls2/genblk1[2].mult/added[2] ), .B(n19733), 
        .Y(n19732) );
  OR2X1 U11860 ( .A(\lamb/scale_ls2/genblk1[2].mult/added[4] ), .B(
        \add_x_64/n1 ), .Y(n18111) );
  NAND3X1 U11861 ( .A(\lamb/scale_ls2/genblk1[2].mult/added[2] ), .B(
        \lamb/scale_ls2/genblk1[2].mult/added[3] ), .C(
        \lamb/scale_ls2/genblk1[2].mult/added[1] ), .Y(n18113) );
  INVX1 U11862 ( .A(n16588), .Y(n18108) );
  AND2X1 U11863 ( .A(n18111), .B(n18108), .Y(n19735) );
  AOI21X1 U11864 ( .A(n18109), .B(n19732), .C(n19735), .Y(
        \lamb/scale_ls3/genblk1[2].mult/logA[0] ) );
  NOR2X1 U11865 ( .A(\lamb/scale_ls2/genblk1[2].mult/added[3] ), .B(n18114), 
        .Y(n18110) );
  NOR3X1 U11866 ( .A(n19733), .B(n19735), .C(n18110), .Y(
        \lamb/scale_ls3/genblk1[2].mult/logA[2] ) );
  NAND3X1 U11867 ( .A(n18111), .B(n17012), .C(n16588), .Y(n18112) );
  OAI21X1 U11868 ( .A(n17012), .B(n16588), .C(n18112), .Y(
        \lamb/scale_ls3/genblk1[2].mult/logA[3] ) );
  INVX1 U11869 ( .A(\lamb/scale_ls2/genblk1[1].mult/added[2] ), .Y(n18150) );
  NOR3X1 U11870 ( .A(\lamb/scale_ls2/genblk1[1].mult/added[3] ), .B(
        \add_x_65/n1 ), .C(\lamb/scale_ls2/genblk1[1].mult/added[4] ), .Y(
        n18115) );
  INVX1 U11871 ( .A(n18115), .Y(n18144) );
  NAND3X1 U11872 ( .A(\lamb/scale_ls2/genblk1[1].mult/added[3] ), .B(
        \add_x_65/n1 ), .C(\lamb/scale_ls2/genblk1[1].mult/added[4] ), .Y(
        n18149) );
  OR2X1 U11873 ( .A(\lamb/scale_ls2/genblk1[1].mult/added[2] ), .B(n16608), 
        .Y(n18131) );
  OAI21X1 U11874 ( .A(n18150), .B(n18144), .C(n18131), .Y(n18139) );
  INVX1 U11875 ( .A(n18139), .Y(n18121) );
  INVX1 U11876 ( .A(\lamb/scale_ls2/genblk1[1].mult/added[1] ), .Y(n18129) );
  NAND2X1 U11877 ( .A(n18129), .B(\lamb/scale_ls2/genblk1[1].mult/added[2] ), 
        .Y(n18127) );
  INVX1 U11878 ( .A(n18127), .Y(n18119) );
  OR2X1 U11879 ( .A(\add_x_65/n1 ), .B(
        \lamb/scale_ls2/genblk1[1].mult/added[4] ), .Y(n18117) );
  AOI21X1 U11880 ( .A(\add_x_65/n1 ), .B(
        \lamb/scale_ls2/genblk1[1].mult/added[4] ), .C(n17013), .Y(n18136) );
  INVX1 U11881 ( .A(n16491), .Y(n18116) );
  AOI21X1 U11882 ( .A(n18116), .B(n16608), .C(n18115), .Y(n18130) );
  INVX1 U11883 ( .A(\lamb/scale_ls2/genblk1[1].mult/added[3] ), .Y(n18145) );
  NAND2X1 U11884 ( .A(\add_x_65/n1 ), .B(
        \lamb/scale_ls2/genblk1[1].mult/added[4] ), .Y(n18125) );
  NAND3X1 U11885 ( .A(n18145), .B(n18125), .C(n18117), .Y(n18138) );
  NAND2X1 U11886 ( .A(n18129), .B(n18138), .Y(n18118) );
  AOI22X1 U11887 ( .A(n18119), .B(n16339), .C(n16912), .D(n18118), .Y(n18120)
         );
  AOI21X1 U11888 ( .A(n18121), .B(n18120), .C(n16746), .Y(n18124) );
  XNOR2X1 U11889 ( .A(n18124), .B(n16322), .Y(n18163) );
  NAND2X1 U11890 ( .A(n18145), .B(n18125), .Y(n18126) );
  AOI22X1 U11891 ( .A(n18129), .B(n17013), .C(n18127), .D(n16425), .Y(n18133)
         );
  NAND2X1 U11892 ( .A(n18131), .B(n16912), .Y(n18132) );
  OAI21X1 U11893 ( .A(n18133), .B(n18132), .C(n18413), .Y(n18135) );
  XNOR2X1 U11894 ( .A(n18135), .B(n16323), .Y(n18160) );
  OR2X1 U11895 ( .A(n18163), .B(n18160), .Y(n18171) );
  INVX1 U11896 ( .A(n16425), .Y(n18137) );
  AOI22X1 U11897 ( .A(\lamb/scale_ls2/genblk1[1].mult/added[2] ), .B(n18137), 
        .C(n16339), .D(n16491), .Y(n18141) );
  INVX1 U11898 ( .A(n18138), .Y(n18147) );
  OAI21X1 U11899 ( .A(n18147), .B(n18139), .C(
        \lamb/scale_ls2/genblk1[1].mult/added[1] ), .Y(n18140) );
  AOI21X1 U11900 ( .A(n18141), .B(n18140), .C(n16746), .Y(n18143) );
  NAND2X1 U11901 ( .A(n17123), .B(n19711), .Y(n18142) );
  HAX1 U11902 ( .A(n16878), .B(n18142), .YS(n18169) );
  OAI21X1 U11903 ( .A(\lamb/scale_ls2/genblk1[1].mult/added[2] ), .B(n18145), 
        .C(n18144), .Y(n18146) );
  AOI22X1 U11904 ( .A(\lamb/scale_ls2/genblk1[1].mult/added[2] ), .B(n18147), 
        .C(\lamb/scale_ls2/genblk1[1].mult/added[1] ), .D(n18146), .Y(n18154)
         );
  OAI21X1 U11905 ( .A(n18150), .B(n16608), .C(n16425), .Y(n18152) );
  AOI21X1 U11906 ( .A(n18154), .B(n16815), .C(n16746), .Y(n18158) );
  NAND2X1 U11907 ( .A(n17123), .B(n18155), .Y(n18157) );
  HAX1 U11908 ( .A(n18158), .B(n18157), .YS(n18164) );
  OR2X1 U11909 ( .A(n18160), .B(n18164), .Y(n18162) );
  OAI21X1 U11910 ( .A(n18173), .B(n18169), .C(n18162), .Y(
        \lamb/scale_ls3/genblk1[1].mult/logA[0] ) );
  INVX1 U11911 ( .A(n18169), .Y(n18159) );
  NAND3X1 U11912 ( .A(n18163), .B(n18169), .C(n18162), .Y(n18161) );
  AND2X1 U11913 ( .A(n18160), .B(n18164), .Y(n18394) );
  AOI21X1 U11914 ( .A(n16341), .B(n18161), .C(n18394), .Y(
        \lamb/scale_ls3/genblk1[1].mult/logA[1] ) );
  INVX1 U11915 ( .A(n18162), .Y(n18168) );
  NAND2X1 U11916 ( .A(n18163), .B(n18169), .Y(n18167) );
  INVX1 U11917 ( .A(n18164), .Y(n18174) );
  OAI21X1 U11918 ( .A(n18167), .B(n18168), .C(n18174), .Y(n18166) );
  AOI22X1 U11919 ( .A(n18168), .B(n18167), .C(n18166), .D(n16341), .Y(
        \lamb/scale_ls3/genblk1[1].mult/logA[2] ) );
  NAND2X1 U11920 ( .A(n17004), .B(n18169), .Y(n18393) );
  OAI21X1 U11921 ( .A(n18171), .B(n18174), .C(n18393), .Y(n18172) );
  AOI21X1 U11922 ( .A(n18174), .B(n18173), .C(n18172), .Y(
        \lamb/scale_ls3/genblk1[1].mult/logA[3] ) );
  NAND2X1 U11923 ( .A(n19770), .B(n18175), .Y(n18176) );
  MUX2X1 U11924 ( .B(n16623), .A(n16392), .S(n18176), .Y(n18177) );
  MUX2X1 U11925 ( .B(n17114), .A(n16617), .S(n16979), .Y(n18182) );
  OAI21X1 U11926 ( .A(n19770), .B(n18182), .C(n16404), .Y(
        \lamb/scale_ls3/genblk1[0].mult/logB[3] ) );
  OAI21X1 U11927 ( .A(n16647), .B(n17102), .C(n18194), .Y(n18185) );
  OAI21X1 U11928 ( .A(n16647), .B(n16610), .C(n17102), .Y(n18435) );
  INVX1 U11929 ( .A(n18435), .Y(n18184) );
  AOI21X1 U11930 ( .A(n18186), .B(n18185), .C(n18184), .Y(
        \lamb/scale_ls3/genblk1[0].mult/logA[1] ) );
  NAND2X1 U11931 ( .A(n17102), .B(n18187), .Y(n18192) );
  INVX1 U11932 ( .A(n16380), .Y(n18188) );
  OAI21X1 U11933 ( .A(n17102), .B(n18188), .C(n18434), .Y(n18189) );
  OAI21X1 U11934 ( .A(n18190), .B(n18192), .C(n18189), .Y(n18191) );
  AOI21X1 U11935 ( .A(n16610), .B(n18192), .C(n18191), .Y(
        \lamb/scale_ls3/genblk1[0].mult/logA[2] ) );
  MUX2X1 U11936 ( .B(n18194), .A(n18434), .S(n16639), .Y(n18196) );
  OAI21X1 U11937 ( .A(n17102), .B(n18196), .C(n16380), .Y(
        \lamb/scale_ls3/genblk1[0].mult/logA[3] ) );
  NAND2X1 U11938 ( .A(n17006), .B(n18202), .Y(n18200) );
  AOI21X1 U11939 ( .A(n19663), .B(n18200), .C(n18199), .Y(
        \lamb/scale_ts2/genblk1[3].mult/logA[1] ) );
  NAND2X1 U11940 ( .A(n18206), .B(n18205), .Y(n18210) );
  AOI21X1 U11941 ( .A(n18202), .B(n19663), .C(n17006), .Y(n18203) );
  AOI21X1 U11942 ( .A(n18210), .B(n18201), .C(n18203), .Y(n18204) );
  OAI21X1 U11943 ( .A(n18206), .B(n18205), .C(n18204), .Y(n18207) );
  INVX1 U11944 ( .A(n18207), .Y(\lamb/scale_ts2/genblk1[3].mult/logA[2] ) );
  INVX1 U11945 ( .A(n18208), .Y(n18211) );
  AOI21X1 U11946 ( .A(n18211), .B(n18210), .C(n18209), .Y(
        \lamb/scale_ts2/genblk1[3].mult/logA[3] ) );
  OAI21X1 U11947 ( .A(n16761), .B(n16663), .C(n16759), .Y(n18215) );
  INVX1 U11948 ( .A(n18213), .Y(n18214) );
  AOI21X1 U11949 ( .A(n16750), .B(n18215), .C(n18214), .Y(
        \lamb/scale_ts2/genblk1[2].mult/logA[1] ) );
  OAI21X1 U11950 ( .A(n18217), .B(n16760), .C(n16761), .Y(n18219) );
  OAI21X1 U11951 ( .A(n16759), .B(n16601), .C(n18219), .Y(n18220) );
  MUX2X1 U11952 ( .B(n18220), .A(n18219), .S(n16650), .Y(
        \lamb/scale_ts2/genblk1[2].mult/logA[2] ) );
  MUX2X1 U11953 ( .B(n16759), .A(n16760), .S(n18221), .Y(n18225) );
  OAI21X1 U11954 ( .A(n18225), .B(n16761), .C(n16601), .Y(
        \lamb/scale_ts2/genblk1[2].mult/logA[3] ) );
  AOI21X1 U11955 ( .A(n18233), .B(n18234), .C(n17024), .Y(n18238) );
  OAI21X1 U11956 ( .A(n16731), .B(n16363), .C(n16574), .Y(
        \lamb/scale_ts2/genblk1[1].mult/logA[0] ) );
  NAND2X1 U11957 ( .A(n18226), .B(n16732), .Y(n18239) );
  AOI21X1 U11958 ( .A(n18228), .B(n16731), .C(n16574), .Y(n18229) );
  AOI21X1 U11959 ( .A(n16731), .B(n16401), .C(n18229), .Y(n18230) );
  INVX1 U11960 ( .A(n18230), .Y(n18231) );
  AOI21X1 U11961 ( .A(n17024), .B(n18239), .C(n18231), .Y(
        \lamb/scale_ts2/genblk1[1].mult/logA[2] ) );
  AND2X1 U11962 ( .A(n18234), .B(n18233), .Y(n18240) );
  NAND2X1 U11963 ( .A(n16401), .B(n16732), .Y(n18237) );
  AOI22X1 U11964 ( .A(n18240), .B(n18239), .C(n16363), .D(n18237), .Y(
        \lamb/scale_ts2/genblk1[1].mult/logA[3] ) );
  INVX1 U11965 ( .A(n19762), .Y(n18242) );
  INVX1 U11966 ( .A(n19759), .Y(n19758) );
  NAND2X1 U11967 ( .A(n19758), .B(n18242), .Y(n18244) );
  OAI21X1 U11968 ( .A(n19765), .B(n18243), .C(n18244), .Y(
        \lamb/scale_ds2/genblk1[3].mult/logA[0] ) );
  NAND2X1 U11969 ( .A(n18245), .B(n18244), .Y(n18248) );
  OAI21X1 U11970 ( .A(n19765), .B(n17062), .C(n18246), .Y(n18247) );
  AOI21X1 U11971 ( .A(n19765), .B(n18248), .C(n18247), .Y(
        \lamb/scale_ds2/genblk1[3].mult/logA[1] ) );
  MUX2X1 U11972 ( .B(n19758), .A(n19759), .S(n17029), .Y(n18249) );
  OAI21X1 U11973 ( .A(n19765), .B(n18249), .C(n17062), .Y(
        \lamb/scale_ds2/genblk1[3].mult/logA[3] ) );
  AOI22X1 U11974 ( .A(n18250), .B(n18254), .C(n18259), .D(n18260), .Y(n18264)
         );
  OAI21X1 U11975 ( .A(n18264), .B(n18258), .C(n18253), .Y(
        \lamb/scale_ds2/genblk1[2].mult/logA[0] ) );
  OAI21X1 U11976 ( .A(n17000), .B(n18254), .C(n18258), .Y(n18251) );
  OAI21X1 U11977 ( .A(n18258), .B(n16345), .C(n18251), .Y(n18252) );
  AOI21X1 U11978 ( .A(n18260), .B(n18261), .C(n18252), .Y(
        \lamb/scale_ds2/genblk1[2].mult/logA[1] ) );
  OR2X1 U11979 ( .A(n18261), .B(n18258), .Y(n18265) );
  OAI21X1 U11980 ( .A(n18262), .B(n18254), .C(n17000), .Y(n18255) );
  OAI21X1 U11981 ( .A(n16863), .B(n16345), .C(n18255), .Y(n18257) );
  AOI21X1 U11982 ( .A(n18261), .B(n18258), .C(n18257), .Y(
        \lamb/scale_ds2/genblk1[2].mult/logA[2] ) );
  NOR2X1 U11983 ( .A(n18260), .B(n18259), .Y(n18266) );
  NAND2X1 U11984 ( .A(n18262), .B(n18261), .Y(n18263) );
  INVX1 U11985 ( .A(n18269), .Y(n18281) );
  OAI21X1 U11986 ( .A(n18274), .B(n18281), .C(n18275), .Y(n18271) );
  NAND3X1 U11987 ( .A(n18278), .B(n18271), .C(n16968), .Y(n18272) );
  AOI21X1 U11988 ( .A(n17075), .B(n18273), .C(n18272), .Y(
        \lamb/scale_ds2/genblk1[1].mult/logA[1] ) );
  OR2X1 U11989 ( .A(n18274), .B(n18287), .Y(n18280) );
  OAI21X1 U11990 ( .A(n17075), .B(n16645), .C(n18275), .Y(n18277) );
  NAND2X1 U11991 ( .A(n17075), .B(n16645), .Y(n18276) );
  NAND3X1 U11992 ( .A(n18278), .B(n18277), .C(n18276), .Y(n18279) );
  AOI21X1 U11993 ( .A(n18281), .B(n18280), .C(n18279), .Y(
        \lamb/scale_ds2/genblk1[1].mult/logA[2] ) );
  INVX1 U11994 ( .A(n18282), .Y(n18285) );
  AOI21X1 U11995 ( .A(n18285), .B(n18284), .C(n16645), .Y(n18291) );
  NAND3X1 U11996 ( .A(n17075), .B(n18287), .C(n17483), .Y(n18290) );
  AOI21X1 U11997 ( .A(n18291), .B(n18290), .C(n16479), .Y(
        \lamb/scale_ds2/genblk1[1].mult/logA[3] ) );
  INVX1 U11998 ( .A(n19725), .Y(n18295) );
  OAI21X1 U11999 ( .A(n16932), .B(n18295), .C(n16381), .Y(n18293) );
  NAND2X1 U12000 ( .A(n16744), .B(n19657), .Y(n19729) );
  AOI22X1 U12001 ( .A(n18295), .B(n16932), .C(n18293), .D(n19729), .Y(
        \lamb/scale_ls2/genblk1[0].mult/logB[2] ) );
  NAND2X1 U12002 ( .A(n16419), .B(n18296), .Y(n18299) );
  AOI21X1 U12003 ( .A(n18300), .B(n18299), .C(n18298), .Y(
        \lamb/scale_ls2/genblk1[0].mult/logA[2] ) );
  AOI21X1 U12004 ( .A(n16661), .B(n18302), .C(n18301), .Y(
        \lamb/scale_ls2/genblk1[0].mult/logA[3] ) );
  NOR2X1 U12005 ( .A(n16653), .B(n17079), .Y(n18304) );
  NOR3X1 U12006 ( .A(n18306), .B(n16376), .C(n18304), .Y(
        \lamb/scale_ts1/genblk1[2].mult/logA[1] ) );
  NAND2X1 U12007 ( .A(n19753), .B(n19751), .Y(n18311) );
  NAND2X1 U12008 ( .A(n19753), .B(n18307), .Y(n18308) );
  MUX2X1 U12009 ( .B(n18309), .A(n16653), .S(n18308), .Y(n18310) );
  AOI21X1 U12010 ( .A(n17079), .B(n18311), .C(n18310), .Y(
        \lamb/scale_ts1/genblk1[2].mult/logA[2] ) );
  INVX1 U12011 ( .A(n19746), .Y(n18316) );
  OAI21X1 U12012 ( .A(n18314), .B(n19743), .C(n19740), .Y(n18313) );
  OAI21X1 U12013 ( .A(n18316), .B(n18315), .C(n18317), .Y(n18312) );
  AOI22X1 U12014 ( .A(n18316), .B(n18313), .C(n19743), .D(n18312), .Y(
        \lamb/scale_ts1/genblk1[1].mult/logA[1] ) );
  MUX2X1 U12015 ( .B(n19740), .A(n18315), .S(n16980), .Y(n18318) );
  OAI21X1 U12016 ( .A(n19743), .B(n18318), .C(n16896), .Y(
        \lamb/scale_ts1/genblk1[1].mult/logA[3] ) );
  NAND3X1 U12017 ( .A(n18323), .B(n18333), .C(n18320), .Y(n18321) );
  AOI22X1 U12018 ( .A(n18322), .B(n18329), .C(n16370), .D(n18321), .Y(
        \lamb/scale_ts1/genblk1[0].mult/logB[1] ) );
  NAND2X1 U12019 ( .A(n18323), .B(n18333), .Y(n18326) );
  OAI21X1 U12020 ( .A(n18326), .B(n18327), .C(n18330), .Y(n18325) );
  AOI22X1 U12021 ( .A(n18327), .B(n18326), .C(n18325), .D(n16370), .Y(
        \lamb/scale_ts1/genblk1[0].mult/logB[2] ) );
  MUX2X1 U12022 ( .B(n18330), .A(n18329), .S(n16982), .Y(n18332) );
  OAI21X1 U12023 ( .A(n18333), .B(n18332), .C(n16482), .Y(
        \lamb/scale_ts1/genblk1[0].mult/logB[3] ) );
  NOR2X1 U12024 ( .A(n18336), .B(n17047), .Y(n18341) );
  INVX1 U12025 ( .A(n18334), .Y(n18335) );
  AOI21X1 U12026 ( .A(n18338), .B(n18337), .C(n17022), .Y(n18340) );
  AOI22X1 U12027 ( .A(n18338), .B(n17047), .C(n18337), .D(n19699), .Y(n18339)
         );
  NOR3X1 U12028 ( .A(n18341), .B(n18340), .C(n18339), .Y(
        \lamb/scale_ds1/genblk1[3].mult/logA[2] ) );
  NOR2X1 U12029 ( .A(n16578), .B(n18341), .Y(n18343) );
  AOI22X1 U12030 ( .A(n18343), .B(n18342), .C(n19699), .D(n17022), .Y(
        \lamb/scale_ds1/genblk1[3].mult/logA[3] ) );
  INVX1 U12031 ( .A(n18346), .Y(n18347) );
  INVX1 U12032 ( .A(n18348), .Y(n18345) );
  AOI22X1 U12033 ( .A(n18348), .B(n18347), .C(n18346), .D(n18345), .Y(n18349)
         );
  INVX1 U12034 ( .A(n18344), .Y(n19724) );
  OAI21X1 U12035 ( .A(n18349), .B(n19724), .C(n16464), .Y(
        \lamb/scale_ds1/genblk1[2].mult/logA[0] ) );
  NAND2X1 U12036 ( .A(n18348), .B(n18347), .Y(n18350) );
  OAI21X1 U12037 ( .A(n19719), .B(n18350), .C(n16883), .Y(n18351) );
  AOI21X1 U12038 ( .A(n19724), .B(n16939), .C(n18351), .Y(
        \lamb/scale_ds1/genblk1[2].mult/logA[3] ) );
  INVX1 U12039 ( .A(n16886), .Y(n18357) );
  OAI21X1 U12040 ( .A(n18356), .B(n18357), .C(n18364), .Y(n18373) );
  NAND2X1 U12041 ( .A(n18353), .B(n18360), .Y(n19737) );
  NAND2X1 U12042 ( .A(n17040), .B(n19737), .Y(n18354) );
  AOI22X1 U12043 ( .A(n18355), .B(n18373), .C(n16702), .D(n18354), .Y(
        \lamb/scale_ds1/genblk1[1].mult/logA[1] ) );
  INVX1 U12044 ( .A(n16398), .Y(n18362) );
  NAND2X1 U12045 ( .A(n18357), .B(n17040), .Y(n18358) );
  MUX2X1 U12046 ( .B(n18362), .A(n16398), .S(n18358), .Y(n18363) );
  NOR2X1 U12047 ( .A(n18360), .B(n16702), .Y(n18370) );
  NAND2X1 U12048 ( .A(n18362), .B(n18361), .Y(n18368) );
  INVX1 U12049 ( .A(n18365), .Y(\lamb/scale_ds1/genblk1[1].mult/logA[2] ) );
  AOI21X1 U12050 ( .A(n18368), .B(n17020), .C(n16702), .Y(n18367) );
  INVX1 U12051 ( .A(n18367), .Y(n19736) );
  AOI22X1 U12052 ( .A(n17020), .B(n18370), .C(n18369), .D(n16787), .Y(n18372)
         );
  OAI21X1 U12053 ( .A(n18373), .B(n19736), .C(n18372), .Y(
        \lamb/scale_ds1/genblk1[1].mult/logA[3] ) );
  OAI21X1 U12054 ( .A(n18376), .B(n18375), .C(n18374), .Y(
        \lamb/scale_ts0/genblk1[1].mult/logA[0] ) );
  OR2X1 U12055 ( .A(n18378), .B(n18377), .Y(n18379) );
  AOI21X1 U12056 ( .A(n17026), .B(n18381), .C(n18379), .Y(
        \lamb/scale_ts0/genblk1[1].mult/logA[1] ) );
  OAI21X1 U12057 ( .A(n18382), .B(n18381), .C(n18380), .Y(n18383) );
  NAND2X1 U12058 ( .A(n18384), .B(n18383), .Y(n18385) );
  AOI22X1 U12059 ( .A(n17026), .B(n16353), .C(n16340), .D(n18385), .Y(
        \lamb/scale_ts0/genblk1[1].mult/logA[2] ) );
  INVX1 U12060 ( .A(\lamb/scale_ls3/genblk1[1].mult/added[1] ), .Y(n18506) );
  NOR2X1 U12061 ( .A(n18506), .B(n16812), .Y(n18541) );
  NAND2X1 U12062 ( .A(\lamb/scale_ls3/genblk1[1].mult/added[3] ), .B(n18455), 
        .Y(n18462) );
  INVX1 U12063 ( .A(\lamb/scale_ls3/genblk1[1].mult/added[3] ), .Y(n18507) );
  INVX1 U12064 ( .A(n16446), .Y(n18390) );
  OAI21X1 U12065 ( .A(n18455), .B(n16326), .C(n18506), .Y(n18537) );
  INVX1 U12066 ( .A(n18537), .Y(n18389) );
  AOI21X1 U12067 ( .A(n18541), .B(n18462), .C(n18389), .Y(n18392) );
  NAND2X1 U12068 ( .A(n18390), .B(n17007), .Y(n18461) );
  INVX1 U12069 ( .A(n18461), .Y(n18457) );
  NAND2X1 U12070 ( .A(n18506), .B(n18457), .Y(n18454) );
  NAND2X1 U12071 ( .A(n18454), .B(n17054), .Y(n18391) );
  AOI22X1 U12072 ( .A(n18392), .B(n17054), .C(
        \lamb/scale_ls3/genblk1[1].mult/added[2] ), .D(n18391), .Y(n18396) );
  INVX1 U12073 ( .A(n18393), .Y(n18395) );
  AOI21X1 U12074 ( .A(n18396), .B(n17021), .C(n18542), .Y(n18411) );
  NOR3X1 U12075 ( .A(\lamb/scale_bs3/genblk1[1].mult/added[3] ), .B(
        \add_x_49/n1 ), .C(\lamb/scale_bs3/genblk1[1].mult/added[4] ), .Y(
        n18523) );
  INVX1 U12076 ( .A(n18523), .Y(n18516) );
  NOR2X1 U12077 ( .A(\add_x_49/n1 ), .B(
        \lamb/scale_bs3/genblk1[1].mult/added[4] ), .Y(n18466) );
  AOI21X1 U12078 ( .A(\lamb/scale_bs3/genblk1[1].mult/added[4] ), .B(
        \add_x_49/n1 ), .C(n18466), .Y(n18515) );
  INVX1 U12079 ( .A(n16440), .Y(n18402) );
  NAND2X1 U12080 ( .A(\lamb/scale_bs3/genblk1[1].mult/added[2] ), .B(n16901), 
        .Y(n18468) );
  INVX1 U12081 ( .A(n18468), .Y(n18400) );
  NAND2X1 U12082 ( .A(\lamb/scale_bs3/genblk1[1].mult/added[1] ), .B(n18516), 
        .Y(n18399) );
  INVX1 U12083 ( .A(\lamb/scale_bs3/genblk1[1].mult/added[2] ), .Y(n18514) );
  AND2X1 U12084 ( .A(\add_x_49/n1 ), .B(
        \lamb/scale_bs3/genblk1[1].mult/added[4] ), .Y(n18397) );
  NAND2X1 U12085 ( .A(n17034), .B(n18399), .Y(n18398) );
  AOI22X1 U12086 ( .A(n18400), .B(n18399), .C(n18514), .D(n18398), .Y(n18409)
         );
  INVX1 U12087 ( .A(\lamb/scale_bs3/genblk1[1].mult/added[1] ), .Y(n18401) );
  INVX1 U12088 ( .A(\lamb/scale_bs3/genblk1[1].mult/added[3] ), .Y(n18467) );
  AOI22X1 U12089 ( .A(\lamb/scale_bs3/genblk1[1].mult/added[3] ), .B(
        \lamb/scale_bs3/genblk1[1].mult/added[1] ), .C(n18401), .D(n18467), 
        .Y(n18472) );
  INVX1 U12090 ( .A(n18472), .Y(n18404) );
  OAI21X1 U12091 ( .A(n18402), .B(\lamb/scale_bs3/genblk1[1].mult/added[1] ), 
        .C(n17034), .Y(n18403) );
  NAND2X1 U12092 ( .A(n18404), .B(n18403), .Y(n18408) );
  NOR2X1 U12093 ( .A(n18406), .B(n18405), .Y(n19782) );
  NAND3X1 U12094 ( .A(n19782), .B(n18407), .C(n19778), .Y(n18970) );
  HAX1 U12095 ( .A(n18411), .B(n16846), .YS(n18823) );
  INVX1 U12096 ( .A(n18823), .Y(n18615) );
  AOI22X1 U12097 ( .A(n18414), .B(n16746), .C(n18156), .D(n18412), .Y(n18415)
         );
  AOI21X1 U12098 ( .A(\add_x_50/n1 ), .B(
        \lamb/scale_bs3/genblk1[0].mult/added[4] ), .C(
        \lamb/scale_bs3/genblk1[0].mult/added[3] ), .Y(n18501) );
  OR2X1 U12099 ( .A(\lamb/scale_bs3/genblk1[0].mult/added[4] ), .B(
        \add_x_50/n1 ), .Y(n18419) );
  NAND2X1 U12100 ( .A(\lamb/scale_bs3/genblk1[0].mult/added[3] ), .B(n18419), 
        .Y(n18421) );
  INVX1 U12101 ( .A(n18421), .Y(n18416) );
  NOR2X1 U12102 ( .A(n16566), .B(n18416), .Y(n18447) );
  AOI22X1 U12103 ( .A(\lamb/scale_bs3/genblk1[0].mult/added[1] ), .B(n18558), 
        .C(\lamb/scale_bs3/genblk1[0].mult/added[2] ), .D(n18447), .Y(n18424)
         );
  INVX1 U12104 ( .A(\lamb/scale_bs3/genblk1[0].mult/added[1] ), .Y(n18561) );
  NAND2X1 U12105 ( .A(\lamb/scale_bs3/genblk1[0].mult/added[4] ), .B(
        \add_x_50/n1 ), .Y(n18417) );
  INVX1 U12106 ( .A(n18417), .Y(n18418) );
  AND2X1 U12107 ( .A(\lamb/scale_bs3/genblk1[0].mult/added[3] ), .B(n18418), 
        .Y(n18448) );
  OR2X1 U12108 ( .A(n18419), .B(\lamb/scale_bs3/genblk1[0].mult/added[3] ), 
        .Y(n18560) );
  NAND3X1 U12109 ( .A(n18560), .B(n18423), .C(
        \lamb/scale_bs3/genblk1[0].mult/added[2] ), .Y(n18420) );
  OAI21X1 U12110 ( .A(\lamb/scale_bs3/genblk1[0].mult/added[2] ), .B(n18448), 
        .C(n18420), .Y(n18503) );
  OAI21X1 U12111 ( .A(n18421), .B(\lamb/scale_bs3/genblk1[0].mult/added[2] ), 
        .C(n18503), .Y(n18422) );
  NAND3X1 U12112 ( .A(n18424), .B(n18423), .C(n16359), .Y(n18425) );
  NAND2X1 U12113 ( .A(n18565), .B(n18425), .Y(n18440) );
  AOI21X1 U12114 ( .A(\lamb/scale_ls3/genblk1[0].mult/added[4] ), .B(
        \add_x_53/n1 ), .C(\lamb/scale_ls3/genblk1[0].mult/added[3] ), .Y(
        n18432) );
  INVX1 U12115 ( .A(n16395), .Y(n18429) );
  NAND2X1 U12116 ( .A(\lamb/scale_ls3/genblk1[0].mult/added[4] ), .B(
        \add_x_53/n1 ), .Y(n18426) );
  OR2X1 U12117 ( .A(\lamb/scale_ls3/genblk1[0].mult/added[4] ), .B(
        \add_x_53/n1 ), .Y(n18430) );
  NAND3X1 U12118 ( .A(\lamb/scale_ls3/genblk1[0].mult/added[3] ), .B(n18426), 
        .C(n18430), .Y(n18441) );
  INVX1 U12119 ( .A(\lamb/scale_ls3/genblk1[0].mult/added[3] ), .Y(n18427) );
  OR2X1 U12120 ( .A(\lamb/scale_ls3/genblk1[0].mult/added[2] ), .B(n16515), 
        .Y(n18496) );
  OAI21X1 U12121 ( .A(n18548), .B(n18496), .C(
        \lamb/scale_ls3/genblk1[0].mult/added[1] ), .Y(n18428) );
  AOI22X1 U12122 ( .A(n18550), .B(n18429), .C(n18441), .D(n18428), .Y(n18438)
         );
  OR2X1 U12123 ( .A(n18430), .B(\lamb/scale_ls3/genblk1[0].mult/added[3] ), 
        .Y(n18491) );
  NAND2X1 U12124 ( .A(\lamb/scale_ls3/genblk1[0].mult/added[3] ), .B(n18430), 
        .Y(n18431) );
  AND2X1 U12125 ( .A(\lamb/scale_ls3/genblk1[0].mult/added[2] ), .B(n16585), 
        .Y(n18437) );
  OAI21X1 U12126 ( .A(n18438), .B(n18437), .C(n18497), .Y(n18439) );
  HAX1 U12127 ( .A(n18440), .B(n18439), .YS(n18710) );
  INVX1 U12128 ( .A(n18710), .Y(n18637) );
  INVX1 U12129 ( .A(n18441), .Y(n18442) );
  INVX1 U12130 ( .A(\lamb/scale_ls3/genblk1[0].mult/added[1] ), .Y(n18493) );
  NAND3X1 U12131 ( .A(n18442), .B(\lamb/scale_ls3/genblk1[0].mult/added[2] ), 
        .C(n18493), .Y(n18498) );
  NAND2X1 U12132 ( .A(n16515), .B(n17044), .Y(n18547) );
  NAND2X1 U12133 ( .A(n16585), .B(\lamb/scale_ls3/genblk1[0].mult/added[1] ), 
        .Y(n18443) );
  NAND3X1 U12134 ( .A(n18498), .B(n18547), .C(n18443), .Y(n18445) );
  AOI21X1 U12135 ( .A(n18491), .B(n17044), .C(n16515), .Y(n18492) );
  OAI21X1 U12136 ( .A(n18445), .B(n18492), .C(n18497), .Y(n18453) );
  OAI21X1 U12137 ( .A(n16335), .B(n18448), .C(n18560), .Y(n18446) );
  INVX1 U12138 ( .A(n18446), .Y(n18500) );
  INVX1 U12139 ( .A(n18447), .Y(n18559) );
  NAND2X1 U12140 ( .A(n18448), .B(n18561), .Y(n18557) );
  OAI21X1 U12141 ( .A(n18559), .B(n18561), .C(n18557), .Y(n18449) );
  INVX1 U12142 ( .A(n18449), .Y(n18450) );
  NAND3X1 U12143 ( .A(n18500), .B(n18450), .C(n18503), .Y(n18451) );
  NAND2X1 U12144 ( .A(n18565), .B(n16795), .Y(n18452) );
  HAX1 U12145 ( .A(n18453), .B(n18452), .YS(n18739) );
  HAX1 U12146 ( .A(n18637), .B(n18739), .YS(n18656) );
  HAX1 U12147 ( .A(n18615), .B(n18656), .YS(n18724) );
  INVX1 U12148 ( .A(n18454), .Y(n18460) );
  NAND3X1 U12149 ( .A(n18507), .B(\lamb/scale_ls3/genblk1[1].mult/added[2] ), 
        .C(n17007), .Y(n18456) );
  NAND2X1 U12150 ( .A(n18456), .B(n17021), .Y(n18538) );
  INVX1 U12151 ( .A(n18538), .Y(n18458) );
  NAND2X1 U12152 ( .A(n18457), .B(n16812), .Y(n18510) );
  AOI22X1 U12153 ( .A(\lamb/scale_ls3/genblk1[1].mult/added[3] ), .B(n18460), 
        .C(\lamb/scale_ls3/genblk1[1].mult/added[1] ), .D(n16840), .Y(n18464)
         );
  AOI21X1 U12154 ( .A(n18464), .B(n18463), .C(n18542), .Y(n18476) );
  OR2X1 U12155 ( .A(n18466), .B(\lamb/scale_bs3/genblk1[1].mult/added[2] ), 
        .Y(n18469) );
  MUX2X1 U12156 ( .B(n18469), .A(n18468), .S(n18467), .Y(n18470) );
  OAI21X1 U12157 ( .A(n18514), .B(n18524), .C(n16903), .Y(n18471) );
  INVX1 U12158 ( .A(n18471), .Y(n18474) );
  AOI21X1 U12159 ( .A(n18474), .B(n16808), .C(n16640), .Y(n18475) );
  HAX1 U12160 ( .A(n18476), .B(n18475), .YS(n18840) );
  INVX1 U12161 ( .A(n18840), .Y(n18822) );
  NAND3X1 U12162 ( .A(\lamb/scale_ls3/genblk1[2].mult/added[3] ), .B(
        \lamb/scale_ls3/genblk1[2].mult/added[4] ), .C(\add_x_51/n1 ), .Y(
        n18577) );
  OR2X1 U12163 ( .A(\lamb/scale_ls3/genblk1[2].mult/added[4] ), .B(
        \add_x_51/n1 ), .Y(n18485) );
  INVX1 U12164 ( .A(n18485), .Y(n18481) );
  INVX1 U12165 ( .A(\lamb/scale_ls3/genblk1[2].mult/added[3] ), .Y(n18574) );
  NAND2X1 U12166 ( .A(n18481), .B(n18574), .Y(n18477) );
  NAND2X1 U12167 ( .A(\lamb/scale_ls3/genblk1[2].mult/added[2] ), .B(n16885), 
        .Y(n18484) );
  INVX1 U12168 ( .A(\lamb/scale_ls3/genblk1[2].mult/added[2] ), .Y(n18488) );
  NAND2X1 U12169 ( .A(\lamb/scale_ls3/genblk1[2].mult/added[1] ), .B(n18488), 
        .Y(n18478) );
  AOI22X1 U12170 ( .A(\lamb/scale_ls3/genblk1[2].mult/added[2] ), .B(n16389), 
        .C(n18484), .D(n18478), .Y(n18587) );
  NAND3X1 U12171 ( .A(\lamb/scale_ls3/genblk1[2].mult/added[4] ), .B(
        \add_x_51/n1 ), .C(n18574), .Y(n18479) );
  OAI21X1 U12172 ( .A(n18485), .B(n18574), .C(n18479), .Y(n18571) );
  NAND2X1 U12173 ( .A(\lamb/scale_ls3/genblk1[2].mult/added[1] ), .B(
        \lamb/scale_ls3/genblk1[2].mult/added[2] ), .Y(n18570) );
  AOI22X1 U12174 ( .A(n18587), .B(n16819), .C(n18571), .D(n18570), .Y(n18483)
         );
  AOI21X1 U12175 ( .A(\add_x_51/n1 ), .B(
        \lamb/scale_ls3/genblk1[2].mult/added[4] ), .C(n18481), .Y(n18580) );
  NAND3X1 U12176 ( .A(n18574), .B(\lamb/scale_ls3/genblk1[2].mult/added[2] ), 
        .C(n16665), .Y(n18482) );
  NAND2X1 U12177 ( .A(n18483), .B(n18482), .Y(n18582) );
  INVX1 U12178 ( .A(n18582), .Y(n18490) );
  INVX1 U12179 ( .A(\lamb/scale_ls3/genblk1[2].mult/added[1] ), .Y(n18575) );
  INVX1 U12180 ( .A(n16389), .Y(n18489) );
  INVX1 U12181 ( .A(n18484), .Y(n18487) );
  INVX1 U12182 ( .A(n16665), .Y(n18586) );
  AOI22X1 U12183 ( .A(\lamb/scale_ls3/genblk1[2].mult/added[3] ), .B(n18586), 
        .C(n18485), .D(n18574), .Y(n18486) );
  AOI22X1 U12184 ( .A(n18489), .B(n18488), .C(n18487), .D(n18486), .Y(n18589)
         );
  HAX1 U12185 ( .A(n18822), .B(n17108), .YS(n18738) );
  INVX1 U12186 ( .A(n18492), .Y(n18495) );
  NAND2X1 U12187 ( .A(n16988), .B(n18493), .Y(n18494) );
  AOI22X1 U12188 ( .A(n18496), .B(n16365), .C(n18495), .D(n18494), .Y(n18499)
         );
  INVX1 U12189 ( .A(n18497), .Y(n18554) );
  AOI21X1 U12190 ( .A(n18499), .B(n18498), .C(n18554), .Y(n18505) );
  OAI21X1 U12191 ( .A(\lamb/scale_bs3/genblk1[0].mult/added[1] ), .B(n16566), 
        .C(n18500), .Y(n18502) );
  AOI21X1 U12192 ( .A(n18503), .B(n18502), .C(n17001), .Y(n18504) );
  HAX1 U12193 ( .A(n16870), .B(n18504), .YS(n18621) );
  NAND3X1 U12194 ( .A(n16810), .B(\lamb/scale_ls3/genblk1[1].mult/added[1] ), 
        .C(\lamb/scale_ls3/genblk1[1].mult/added[2] ), .Y(n18511) );
  OAI21X1 U12195 ( .A(n16446), .B(n18507), .C(n18506), .Y(n18509) );
  NAND3X1 U12196 ( .A(n18511), .B(n18510), .C(n18509), .Y(n18512) );
  AOI21X1 U12197 ( .A(n17054), .B(n18512), .C(n18542), .Y(n18522) );
  NAND2X1 U12198 ( .A(\lamb/scale_bs3/genblk1[1].mult/added[2] ), .B(
        \lamb/scale_bs3/genblk1[1].mult/added[1] ), .Y(n18520) );
  OAI21X1 U12199 ( .A(n18514), .B(n18526), .C(n18524), .Y(n18529) );
  INVX1 U12200 ( .A(n18529), .Y(n18518) );
  AOI21X1 U12201 ( .A(n16440), .B(\lamb/scale_bs3/genblk1[1].mult/added[3] ), 
        .C(\lamb/scale_bs3/genblk1[1].mult/added[1] ), .Y(n18517) );
  OAI21X1 U12202 ( .A(n18518), .B(n18517), .C(n18516), .Y(n18519) );
  AOI21X1 U12203 ( .A(n18526), .B(n18520), .C(n18519), .Y(n18530) );
  OR2X1 U12204 ( .A(n18530), .B(n16640), .Y(n18521) );
  HAX1 U12205 ( .A(n18522), .B(n18521), .YS(n19261) );
  AOI21X1 U12206 ( .A(n18523), .B(\lamb/scale_bs3/genblk1[1].mult/added[1] ), 
        .C(\lamb/scale_bs3/genblk1[1].mult/added[2] ), .Y(n18525) );
  AOI22X1 U12207 ( .A(\lamb/scale_bs3/genblk1[1].mult/added[1] ), .B(
        \lamb/scale_bs3/genblk1[1].mult/added[2] ), .C(n18525), .D(n18524), 
        .Y(n18528) );
  NAND2X1 U12208 ( .A(\lamb/scale_bs3/genblk1[1].mult/added[2] ), .B(n17034), 
        .Y(n18527) );
  AOI22X1 U12209 ( .A(n18530), .B(n18529), .C(n18528), .D(n18527), .Y(n18533)
         );
  AOI21X1 U12210 ( .A(n18533), .B(n16903), .C(n16640), .Y(n18545) );
  AOI22X1 U12211 ( .A(\lamb/scale_ls3/genblk1[1].mult/added[1] ), .B(n16326), 
        .C(n18535), .D(n17021), .Y(n18540) );
  NAND2X1 U12212 ( .A(n18538), .B(n18537), .Y(n18539) );
  OAI21X1 U12213 ( .A(n18541), .B(n18540), .C(n18539), .Y(n18543) );
  NAND2X1 U12214 ( .A(n18543), .B(n16884), .Y(n18544) );
  HAX1 U12215 ( .A(n18545), .B(n18544), .YS(n18821) );
  XNOR2X1 U12216 ( .A(n19261), .B(n18821), .Y(n18838) );
  HAX1 U12217 ( .A(n18621), .B(n18838), .YS(n18633) );
  INVX1 U12218 ( .A(n18633), .Y(n18546) );
  HAX1 U12219 ( .A(n18738), .B(n18546), .YS(n18696) );
  INVX1 U12220 ( .A(n18821), .Y(n18598) );
  NAND2X1 U12221 ( .A(n18598), .B(n18840), .Y(n18825) );
  NAND2X1 U12222 ( .A(n16988), .B(n18547), .Y(n18549) );
  AOI22X1 U12223 ( .A(n16585), .B(n17044), .C(
        \lamb/scale_ls3/genblk1[0].mult/added[2] ), .D(n18549), .Y(n18556) );
  NAND3X1 U12224 ( .A(\lamb/scale_ls3/genblk1[0].mult/added[1] ), .B(n16926), 
        .C(n16365), .Y(n18555) );
  AOI21X1 U12225 ( .A(n18556), .B(n18555), .C(n18554), .Y(n18569) );
  NAND2X1 U12226 ( .A(n16887), .B(n18557), .Y(n18564) );
  OAI21X1 U12227 ( .A(n18561), .B(n18560), .C(n18559), .Y(n18562) );
  AOI22X1 U12228 ( .A(\lamb/scale_bs3/genblk1[0].mult/added[2] ), .B(n18564), 
        .C(n16335), .D(n18562), .Y(n18567) );
  AOI21X1 U12229 ( .A(n18567), .B(n16359), .C(n17001), .Y(n18568) );
  HAX1 U12230 ( .A(n18569), .B(n18568), .YS(n18607) );
  XNOR2X1 U12231 ( .A(n18621), .B(n18607), .Y(n18631) );
  HAX1 U12232 ( .A(n18615), .B(n18631), .YS(n18667) );
  INVX1 U12233 ( .A(n18570), .Y(n18585) );
  AOI22X1 U12234 ( .A(\lamb/scale_ls3/genblk1[2].mult/added[3] ), .B(n18585), 
        .C(n18575), .D(n18574), .Y(n18572) );
  AOI22X1 U12235 ( .A(n16665), .B(n18572), .C(
        \lamb/scale_ls3/genblk1[2].mult/added[2] ), .D(n18571), .Y(n18584) );
  HAX1 U12236 ( .A(n18667), .B(n17116), .YS(n18657) );
  AND2X1 U12237 ( .A(n18575), .B(n18574), .Y(n18579) );
  NAND2X1 U12238 ( .A(\lamb/scale_ls3/genblk1[2].mult/added[2] ), .B(n16389), 
        .Y(n18578) );
  AOI22X1 U12239 ( .A(n16665), .B(n18579), .C(n18576), .D(n18578), .Y(n18581)
         );
  HAX1 U12240 ( .A(n18607), .B(n17115), .YS(n18599) );
  XNOR2X1 U12241 ( .A(n18615), .B(n18838), .Y(n18630) );
  HAX1 U12242 ( .A(n18599), .B(n18630), .YS(n18593) );
  INVX1 U12243 ( .A(n18838), .Y(n18670) );
  OAI21X1 U12244 ( .A(n18582), .B(n17115), .C(n16533), .Y(n18583) );
  OAI21X1 U12245 ( .A(n18585), .B(n16533), .C(n18583), .Y(n18590) );
  XNOR2X1 U12246 ( .A(n18607), .B(n16764), .Y(n18729) );
  XNOR2X1 U12247 ( .A(n18822), .B(n18710), .Y(n18746) );
  FAX1 U12248 ( .A(n18670), .B(n18729), .C(n18746), .YS(n18591) );
  OAI21X1 U12249 ( .A(n18739), .B(n18593), .C(n18591), .Y(n18592) );
  AOI21X1 U12250 ( .A(n18739), .B(n18593), .C(n18592), .Y(n18594) );
  OAI21X1 U12251 ( .A(n17072), .B(n18657), .C(n18594), .Y(n18595) );
  AOI21X1 U12252 ( .A(n17072), .B(n18657), .C(n18595), .Y(n18596) );
  OAI21X1 U12253 ( .A(n18724), .B(n18696), .C(n18596), .Y(n18597) );
  AOI21X1 U12254 ( .A(n18724), .B(n18696), .C(n18597), .Y(n18954) );
  HAX1 U12255 ( .A(n19261), .B(n17072), .YS(n18688) );
  HAX1 U12256 ( .A(n18656), .B(n17116), .YS(n18644) );
  HAX1 U12257 ( .A(n18607), .B(n18598), .YS(n18737) );
  XNOR2X1 U12258 ( .A(n18615), .B(n18710), .Y(n18708) );
  HAX1 U12259 ( .A(n18738), .B(n18708), .YS(n18679) );
  INVX1 U12260 ( .A(n18599), .Y(n18709) );
  HAX1 U12261 ( .A(n18621), .B(n18709), .YS(n18664) );
  XNOR2X1 U12262 ( .A(n18615), .B(n18822), .Y(n18837) );
  HAX1 U12263 ( .A(n18838), .B(n18837), .YS(n18601) );
  HAX1 U12264 ( .A(n16764), .B(n18837), .YS(n18632) );
  HAX1 U12265 ( .A(n18621), .B(n18632), .YS(n18606) );
  OAI21X1 U12266 ( .A(n18664), .B(n18601), .C(n18606), .Y(n18600) );
  AOI21X1 U12267 ( .A(n18664), .B(n18601), .C(n18600), .Y(n18602) );
  OAI21X1 U12268 ( .A(n18737), .B(n18679), .C(n16789), .Y(n18603) );
  AOI21X1 U12269 ( .A(n18737), .B(n18679), .C(n18603), .Y(n18604) );
  OAI21X1 U12270 ( .A(n18688), .B(n18644), .C(n18604), .Y(n18605) );
  AOI21X1 U12271 ( .A(n18688), .B(n18644), .C(n18605), .Y(n18763) );
  INVX1 U12272 ( .A(n18763), .Y(n18908) );
  INVX1 U12273 ( .A(n18606), .Y(n18681) );
  XNOR2X1 U12274 ( .A(n18821), .B(n18710), .Y(n18736) );
  HAX1 U12275 ( .A(n18739), .B(n18736), .YS(n18693) );
  INVX1 U12276 ( .A(n18693), .Y(n18697) );
  HAX1 U12277 ( .A(n18739), .B(n18670), .YS(n18678) );
  XNOR2X1 U12278 ( .A(n18607), .B(n17116), .Y(n18707) );
  XNOR2X1 U12279 ( .A(n18837), .B(n18707), .Y(n18694) );
  NAND2X1 U12280 ( .A(n18823), .B(n19261), .Y(n18824) );
  NAND2X1 U12281 ( .A(n16996), .B(n18615), .Y(n18819) );
  HAX1 U12282 ( .A(n18656), .B(n18709), .YS(n18610) );
  INVX1 U12283 ( .A(n18736), .Y(n18727) );
  HAX1 U12284 ( .A(n18621), .B(n17108), .YS(n18669) );
  HAX1 U12285 ( .A(n18727), .B(n18669), .YS(n18608) );
  MUX2X1 U12286 ( .B(n18610), .A(n18833), .S(n18608), .Y(n18609) );
  AOI21X1 U12287 ( .A(n18833), .B(n18610), .C(n18609), .Y(n18611) );
  AOI21X1 U12288 ( .A(n18681), .B(n18697), .C(n16798), .Y(n18614) );
  OAI21X1 U12289 ( .A(n18681), .B(n18697), .C(n18614), .Y(n19264) );
  INVX1 U12290 ( .A(n19264), .Y(n18905) );
  HAX1 U12291 ( .A(n18737), .B(n17108), .YS(n18719) );
  HAX1 U12292 ( .A(n16996), .B(n16764), .YS(n18645) );
  INVX1 U12293 ( .A(n18645), .Y(n18622) );
  INVX1 U12294 ( .A(n18746), .Y(n18618) );
  HAX1 U12295 ( .A(n18621), .B(n17115), .YS(n18649) );
  INVX1 U12296 ( .A(n18649), .Y(n18701) );
  XNOR2X1 U12297 ( .A(n18615), .B(n18701), .Y(n18735) );
  INVX1 U12298 ( .A(n18735), .Y(n18616) );
  AOI21X1 U12299 ( .A(n17116), .B(n18618), .C(n18616), .Y(n18617) );
  OAI21X1 U12300 ( .A(n17116), .B(n18618), .C(n18617), .Y(n18619) );
  AOI21X1 U12301 ( .A(n18739), .B(n18622), .C(n18619), .Y(n18620) );
  OAI21X1 U12302 ( .A(n18739), .B(n18622), .C(n18620), .Y(n18629) );
  HAX1 U12303 ( .A(n18621), .B(n17116), .YS(n18726) );
  HAX1 U12304 ( .A(n19261), .B(n18739), .YS(n18728) );
  HAX1 U12305 ( .A(n18726), .B(n18728), .YS(n18745) );
  HAX1 U12306 ( .A(n18667), .B(n18622), .YS(n18623) );
  MUX2X1 U12307 ( .B(n18739), .A(n18738), .S(n18623), .Y(n18624) );
  AOI21X1 U12308 ( .A(n18738), .B(n18739), .C(n18624), .Y(n18625) );
  NAND2X1 U12309 ( .A(n18745), .B(n18625), .Y(n18626) );
  AOI21X1 U12310 ( .A(n17115), .B(n18727), .C(n18626), .Y(n18627) );
  OAI21X1 U12311 ( .A(n17115), .B(n18727), .C(n18627), .Y(n18628) );
  OAI21X1 U12312 ( .A(n18719), .B(n18629), .C(n18628), .Y(n18912) );
  INVX1 U12313 ( .A(n18912), .Y(n18906) );
  HAX1 U12314 ( .A(n18630), .B(n18707), .YS(n18643) );
  HAX1 U12315 ( .A(n19261), .B(n18631), .YS(n18704) );
  INVX1 U12316 ( .A(n18704), .Y(n18668) );
  HAX1 U12317 ( .A(n18668), .B(n18656), .YS(n18658) );
  INVX1 U12318 ( .A(n18658), .Y(n18640) );
  HAX1 U12319 ( .A(n18631), .B(n17066), .YS(n18721) );
  XNOR2X1 U12320 ( .A(n18721), .B(n17108), .Y(n18636) );
  HAX1 U12321 ( .A(n18633), .B(n18632), .YS(n18634) );
  MUX2X1 U12322 ( .B(n18636), .A(n18637), .S(n18634), .Y(n18635) );
  OAI21X1 U12323 ( .A(n18637), .B(n18636), .C(n18635), .Y(n18638) );
  AOI21X1 U12324 ( .A(n17115), .B(n18640), .C(n18638), .Y(n18639) );
  OAI21X1 U12325 ( .A(n17115), .B(n18640), .C(n18639), .Y(n18641) );
  AOI21X1 U12326 ( .A(n18656), .B(n18643), .C(n18641), .Y(n18642) );
  OAI21X1 U12327 ( .A(n18656), .B(n18643), .C(n18642), .Y(n18766) );
  INVX1 U12328 ( .A(n18644), .Y(n18648) );
  HAX1 U12329 ( .A(n18727), .B(n18645), .YS(n18690) );
  HAX1 U12330 ( .A(n18667), .B(n18690), .YS(n18646) );
  OAI21X1 U12331 ( .A(n18648), .B(n18721), .C(n18646), .Y(n18647) );
  AOI21X1 U12332 ( .A(n18648), .B(n18721), .C(n18647), .Y(n18654) );
  HAX1 U12333 ( .A(n18668), .B(n17108), .YS(n18652) );
  HAX1 U12334 ( .A(n18822), .B(n18649), .YS(n18650) );
  MUX2X1 U12335 ( .B(n18739), .A(n18652), .S(n18650), .Y(n18651) );
  AOI21X1 U12336 ( .A(n18652), .B(n18739), .C(n18651), .Y(n18653) );
  NAND2X1 U12337 ( .A(n18654), .B(n18653), .Y(n18754) );
  NAND2X1 U12338 ( .A(n18766), .B(n18754), .Y(n18755) );
  INVX1 U12339 ( .A(n18755), .Y(n18768) );
  HAX1 U12340 ( .A(n18656), .B(n17072), .YS(n18700) );
  INVX1 U12341 ( .A(n18657), .Y(n18661) );
  FAX1 U12342 ( .A(n18837), .B(n18658), .C(n17108), .YS(n18659) );
  OAI21X1 U12343 ( .A(n18736), .B(n18661), .C(n18659), .Y(n18660) );
  AOI21X1 U12344 ( .A(n18736), .B(n18661), .C(n18660), .Y(n18662) );
  OAI21X1 U12345 ( .A(n18664), .B(n18678), .C(n16792), .Y(n18663) );
  AOI21X1 U12346 ( .A(n18664), .B(n18678), .C(n18663), .Y(n18665) );
  OAI21X1 U12347 ( .A(n18729), .B(n18700), .C(n18665), .Y(n18666) );
  AOI21X1 U12348 ( .A(n18729), .B(n18700), .C(n18666), .Y(n18815) );
  INVX1 U12349 ( .A(n16748), .Y(n18791) );
  XNOR2X1 U12350 ( .A(n18667), .B(n16764), .Y(n18740) );
  XNOR2X1 U12351 ( .A(n18837), .B(n17115), .Y(n18689) );
  FAX1 U12352 ( .A(n18837), .B(n17116), .C(n18668), .YS(n18671) );
  NOR3X1 U12353 ( .A(n18689), .B(n18671), .C(n18739), .Y(n18675) );
  HAX1 U12354 ( .A(n18670), .B(n18669), .YS(n18674) );
  NAND3X1 U12355 ( .A(n18689), .B(n18671), .C(n18739), .Y(n18672) );
  OAI21X1 U12356 ( .A(n18675), .B(n18674), .C(n16790), .Y(n18676) );
  AOI21X1 U12357 ( .A(n18693), .B(n18740), .C(n18676), .Y(n18677) );
  OAI21X1 U12358 ( .A(n18693), .B(n18740), .C(n18677), .Y(n18940) );
  AND2X1 U12359 ( .A(n18791), .B(n18940), .Y(n18915) );
  INVX1 U12360 ( .A(n18678), .Y(n18684) );
  OAI21X1 U12361 ( .A(n18681), .B(n18728), .C(n18679), .Y(n18680) );
  AOI21X1 U12362 ( .A(n18681), .B(n18728), .C(n18680), .Y(n18682) );
  OAI21X1 U12363 ( .A(n17116), .B(n18684), .C(n18682), .Y(n18683) );
  AOI21X1 U12364 ( .A(n17116), .B(n18684), .C(n18683), .Y(n18686) );
  OAI21X1 U12365 ( .A(n18709), .B(n18688), .C(n18686), .Y(n18687) );
  AOI21X1 U12366 ( .A(n18709), .B(n18688), .C(n18687), .Y(n18764) );
  INVX1 U12367 ( .A(n18764), .Y(n18938) );
  INVX1 U12368 ( .A(n18689), .Y(n18692) );
  OAI21X1 U12369 ( .A(n18693), .B(n18692), .C(n18690), .Y(n18691) );
  AOI21X1 U12370 ( .A(n18693), .B(n18692), .C(n18691), .Y(n18695) );
  NAND3X1 U12371 ( .A(n18696), .B(n18695), .C(n18694), .Y(n18941) );
  INVX1 U12372 ( .A(n16512), .Y(n19547) );
  HAX1 U12373 ( .A(n16764), .B(n18697), .YS(n18698) );
  OAI21X1 U12374 ( .A(n18701), .B(n18700), .C(n18698), .Y(n18699) );
  AOI21X1 U12375 ( .A(n18701), .B(n18700), .C(n18699), .Y(n18702) );
  OAI21X1 U12376 ( .A(n18738), .B(n18704), .C(n18702), .Y(n18703) );
  AOI21X1 U12377 ( .A(n18738), .B(n18704), .C(n18703), .Y(n18705) );
  OAI21X1 U12378 ( .A(n18708), .B(n18707), .C(n18705), .Y(n18706) );
  AOI21X1 U12379 ( .A(n18708), .B(n18707), .C(n18706), .Y(n18928) );
  INVX1 U12380 ( .A(n16379), .Y(n18898) );
  INVX1 U12381 ( .A(n18724), .Y(n18718) );
  HAX1 U12382 ( .A(n18821), .B(n18726), .YS(n18714) );
  FAX1 U12383 ( .A(n16996), .B(n18710), .C(n18709), .YS(n18711) );
  MUX2X1 U12384 ( .B(n18840), .A(n18729), .S(n18711), .Y(n18712) );
  AOI21X1 U12385 ( .A(n18729), .B(n18840), .C(n18712), .Y(n18713) );
  NAND2X1 U12386 ( .A(n18714), .B(n18713), .Y(n18715) );
  AOI21X1 U12387 ( .A(n18718), .B(n17108), .C(n18715), .Y(n18716) );
  OAI21X1 U12388 ( .A(n18718), .B(n17108), .C(n18716), .Y(n18808) );
  NAND2X1 U12389 ( .A(n18898), .B(n18808), .Y(n18747) );
  INVX1 U12390 ( .A(n18719), .Y(n18725) );
  FAX1 U12391 ( .A(n18746), .B(n18721), .C(n17115), .YS(n18722) );
  OAI21X1 U12392 ( .A(n18725), .B(n18724), .C(n18722), .Y(n18723) );
  AOI21X1 U12393 ( .A(n18725), .B(n18724), .C(n18723), .Y(n18734) );
  HAX1 U12394 ( .A(n18727), .B(n18726), .YS(n18732) );
  XNOR2X1 U12395 ( .A(n18729), .B(n18728), .Y(n18730) );
  MUX2X1 U12396 ( .B(n18840), .A(n18732), .S(n18730), .Y(n18731) );
  AOI21X1 U12397 ( .A(n18732), .B(n18840), .C(n18731), .Y(n18733) );
  HAX1 U12398 ( .A(n18736), .B(n18735), .YS(n18742) );
  FAX1 U12399 ( .A(n18739), .B(n18738), .C(n18737), .YS(n18741) );
  NAND3X1 U12400 ( .A(n18742), .B(n18741), .C(n18740), .Y(n18743) );
  AOI21X1 U12401 ( .A(n18746), .B(n18745), .C(n16797), .Y(n18744) );
  OAI21X1 U12402 ( .A(n18746), .B(n18745), .C(n18744), .Y(n18757) );
  INVX1 U12403 ( .A(n18816), .Y(n18812) );
  NOR3X1 U12404 ( .A(n16921), .B(n16576), .C(n16338), .Y(n18751) );
  NAND2X1 U12405 ( .A(n18752), .B(n18751), .Y(n18753) );
  NAND3X1 U12406 ( .A(n19623), .B(n18812), .C(n18753), .Y(valid) );
  NAND2X1 U12407 ( .A(n16660), .B(n18766), .Y(n18760) );
  NAND2X1 U12408 ( .A(n18905), .B(n18755), .Y(n18776) );
  NAND2X1 U12409 ( .A(n17107), .B(n16644), .Y(n18759) );
  NAND2X1 U12410 ( .A(n18759), .B(n16563), .Y(n18756) );
  OR2X1 U12411 ( .A(n18945), .B(n16416), .Y(n18781) );
  INVX1 U12412 ( .A(n18757), .Y(n18927) );
  NAND2X1 U12413 ( .A(n18915), .B(n16914), .Y(n18926) );
  NAND3X1 U12414 ( .A(n17078), .B(n18926), .C(n18945), .Y(n18780) );
  NAND3X1 U12415 ( .A(n18917), .B(n18781), .C(n18780), .Y(n18758) );
  AOI21X1 U12416 ( .A(n17101), .B(n18758), .C(n16506), .Y(n18762) );
  NAND3X1 U12417 ( .A(n16413), .B(n18760), .C(n18759), .Y(n18761) );
  NOR2X1 U12418 ( .A(n18784), .B(n16473), .Y(n18792) );
  OAI21X1 U12419 ( .A(n18792), .B(n16748), .C(n18934), .Y(n18765) );
  NAND2X1 U12420 ( .A(n16723), .B(n18765), .Y(n18773) );
  NAND2X1 U12421 ( .A(n16762), .B(n18773), .Y(n18775) );
  INVX1 U12422 ( .A(n18775), .Y(n18767) );
  OAI21X1 U12423 ( .A(n16657), .B(n18767), .C(n18766), .Y(n19448) );
  NAND2X1 U12424 ( .A(n18768), .B(n19264), .Y(n19259) );
  OAI21X1 U12425 ( .A(n17078), .B(n16748), .C(n16379), .Y(n18896) );
  INVX1 U12426 ( .A(n18896), .Y(n18772) );
  INVX1 U12427 ( .A(n16473), .Y(n18770) );
  AOI22X1 U12428 ( .A(n18791), .B(n18944), .C(n16626), .D(n18770), .Y(n18771)
         );
  NOR3X1 U12429 ( .A(n18772), .B(n17107), .C(n18771), .Y(n18794) );
  OR2X1 U12430 ( .A(n18940), .B(n18945), .Y(n18929) );
  AOI22X1 U12431 ( .A(n18794), .B(n18929), .C(n17107), .D(n18773), .Y(n18774)
         );
  NAND2X1 U12432 ( .A(n16825), .B(n18774), .Y(n18778) );
  NAND3X1 U12433 ( .A(n18778), .B(n18777), .C(n18906), .Y(n18779) );
  OAI21X1 U12434 ( .A(n18906), .B(n19448), .C(n18779), .Y(n19620) );
  INVX1 U12435 ( .A(n18780), .Y(n18805) );
  INVX1 U12436 ( .A(n18781), .Y(n18782) );
  NAND3X1 U12437 ( .A(n19256), .B(n18782), .C(n16583), .Y(n18803) );
  OR2X1 U12438 ( .A(n16644), .B(n16620), .Y(n19523) );
  INVX1 U12439 ( .A(n19523), .Y(n18786) );
  MUX2X1 U12440 ( .B(n16763), .A(n18952), .S(n18786), .Y(n18813) );
  NAND2X1 U12441 ( .A(n18905), .B(n17074), .Y(n18799) );
  NAND3X1 U12442 ( .A(n19268), .B(n18813), .C(n18799), .Y(n18802) );
  OAI21X1 U12443 ( .A(n16735), .B(n17107), .C(n16625), .Y(n18785) );
  AOI21X1 U12444 ( .A(n16658), .B(n17107), .C(n18785), .Y(n18790) );
  AOI21X1 U12445 ( .A(n18938), .B(n16625), .C(n17107), .Y(n19260) );
  AOI22X1 U12446 ( .A(n19260), .B(n19523), .C(n16644), .D(n16506), .Y(n18789)
         );
  OAI21X1 U12447 ( .A(n18790), .B(n16952), .C(n18789), .Y(n18857) );
  AND2X1 U12448 ( .A(n18937), .B(n18917), .Y(n19549) );
  OAI21X1 U12449 ( .A(n18792), .B(n16940), .C(n16723), .Y(n18793) );
  INVX1 U12450 ( .A(n18793), .Y(n18796) );
  AOI21X1 U12451 ( .A(n18908), .B(n18796), .C(n16763), .Y(n19270) );
  AOI22X1 U12452 ( .A(n19549), .B(n18794), .C(n19523), .D(n17059), .Y(n18800)
         );
  NOR2X1 U12453 ( .A(n19523), .B(n18952), .Y(n18797) );
  NAND3X1 U12454 ( .A(n18797), .B(n18796), .C(n16563), .Y(n18798) );
  OR2X1 U12455 ( .A(n18857), .B(n16724), .Y(n18801) );
  NAND3X1 U12456 ( .A(n18803), .B(n18802), .C(n18801), .Y(n18804) );
  AOI21X1 U12457 ( .A(n18937), .B(n18805), .C(n18804), .Y(n18848) );
  AND2X1 U12458 ( .A(n18917), .B(n18929), .Y(n18949) );
  OAI21X1 U12459 ( .A(n18808), .B(n18898), .C(n16416), .Y(n18810) );
  NAND3X1 U12460 ( .A(n18808), .B(n18898), .C(n16914), .Y(n18809) );
  NAND2X1 U12461 ( .A(n18810), .B(n18809), .Y(n18811) );
  OAI21X1 U12462 ( .A(n16748), .B(n18812), .C(n18944), .Y(n19258) );
  AOI22X1 U12463 ( .A(n18937), .B(n16820), .C(n18813), .D(n19258), .Y(n18818)
         );
  NAND2X1 U12464 ( .A(n17074), .B(n16657), .Y(n18957) );
  NAND3X1 U12465 ( .A(n19570), .B(n18816), .C(n16930), .Y(n18817) );
  MUX2X1 U12466 ( .B(n17066), .A(n18819), .S(n18821), .Y(n18820) );
  OAI21X1 U12467 ( .A(n18822), .B(n18820), .C(n18824), .Y(n19267) );
  NOR2X1 U12468 ( .A(n19261), .B(n18821), .Y(n18832) );
  NAND2X1 U12469 ( .A(n18823), .B(n18822), .Y(n18827) );
  INVX1 U12470 ( .A(n18824), .Y(n18826) );
  AOI22X1 U12471 ( .A(n18832), .B(n18827), .C(n18826), .D(n18825), .Y(n18829)
         );
  AND2X1 U12472 ( .A(n18829), .B(n16551), .Y(n19272) );
  OR2X1 U12473 ( .A(n18830), .B(n19272), .Y(n18835) );
  NAND3X1 U12474 ( .A(n19262), .B(n18835), .C(n16900), .Y(n18831) );
  HAX1 U12475 ( .A(n16587), .B(n18831), .YS(n18886) );
  INVX1 U12476 ( .A(n18886), .Y(n18884) );
  NAND2X1 U12477 ( .A(n17046), .B(n19262), .Y(n18844) );
  AOI21X1 U12478 ( .A(n18840), .B(n17066), .C(n18832), .Y(n19282) );
  OAI21X1 U12479 ( .A(n16587), .B(n18834), .C(n18835), .Y(n18841) );
  NOR2X1 U12480 ( .A(n18838), .B(n18837), .Y(n18839) );
  AOI21X1 U12481 ( .A(n18840), .B(n16996), .C(n18839), .Y(n19275) );
  NOR2X1 U12482 ( .A(n18841), .B(n17043), .Y(n18851) );
  NAND2X1 U12483 ( .A(n17043), .B(n18841), .Y(n18853) );
  OAI21X1 U12484 ( .A(n18851), .B(n16724), .C(n18853), .Y(n18842) );
  NAND2X1 U12485 ( .A(n16648), .B(n18842), .Y(n18847) );
  OR2X1 U12486 ( .A(n18842), .B(n16648), .Y(n18846) );
  NAND2X1 U12487 ( .A(n18847), .B(n18846), .Y(n18843) );
  MUX2X1 U12488 ( .B(n18844), .A(n17046), .S(n18843), .Y(n18888) );
  INVX1 U12489 ( .A(n18888), .Y(n18874) );
  HAX1 U12490 ( .A(n16470), .B(n16612), .YS(n18882) );
  AND2X1 U12491 ( .A(n19262), .B(n18846), .Y(n18850) );
  NAND2X1 U12492 ( .A(n17046), .B(n18847), .Y(n18849) );
  OR2X1 U12493 ( .A(n18882), .B(n16641), .Y(n18891) );
  INVX1 U12494 ( .A(n18851), .Y(n18852) );
  NAND3X1 U12495 ( .A(n19262), .B(n18853), .C(n18852), .Y(n18854) );
  HAX1 U12496 ( .A(n16724), .B(n18854), .YS(n18876) );
  INVX1 U12497 ( .A(n18876), .Y(n18866) );
  NAND2X1 U12498 ( .A(n18856), .B(n18888), .Y(n18855) );
  OAI21X1 U12499 ( .A(n18886), .B(n18866), .C(n18855), .Y(n18889) );
  AND2X1 U12500 ( .A(n18874), .B(n18891), .Y(n18885) );
  MUX2X1 U12501 ( .B(n18866), .A(n16898), .S(n18885), .Y(n18861) );
  INVX1 U12502 ( .A(n18857), .Y(n18860) );
  NAND2X1 U12503 ( .A(n16618), .B(n19261), .Y(n18858) );
  OAI21X1 U12504 ( .A(n18860), .B(n16554), .C(n18858), .Y(n18865) );
  AOI21X1 U12505 ( .A(n18861), .B(n17092), .C(n18865), .Y(n18862) );
  OAI21X1 U12506 ( .A(n17092), .B(n18889), .C(n18862), .Y(n18863) );
  INVX1 U12507 ( .A(n18863), .Y(n18864) );
  OAI21X1 U12508 ( .A(n16928), .B(n18891), .C(n18864), .Y(n19209) );
  INVX1 U12509 ( .A(n19209), .Y(n19215) );
  INVX1 U12510 ( .A(n18865), .Y(n18895) );
  INVX1 U12511 ( .A(n18882), .Y(n18887) );
  AOI21X1 U12512 ( .A(n18876), .B(n18886), .C(n16641), .Y(n18870) );
  NAND2X1 U12513 ( .A(n16641), .B(n18866), .Y(n18881) );
  NAND3X1 U12514 ( .A(n16928), .B(n18881), .C(n18887), .Y(n18869) );
  OAI21X1 U12515 ( .A(n18887), .B(n18870), .C(n18869), .Y(n18873) );
  NOR2X1 U12516 ( .A(n18888), .B(n17092), .Y(n18871) );
  NAND2X1 U12517 ( .A(n18886), .B(n18871), .Y(n18872) );
  NAND3X1 U12518 ( .A(n18895), .B(n18873), .C(n18872), .Y(n19204) );
  INVX1 U12519 ( .A(n19204), .Y(n19210) );
  MUX2X1 U12520 ( .B(n18876), .A(n17092), .S(n18874), .Y(n18879) );
  MUX2X1 U12521 ( .B(n18888), .A(n18876), .S(n17092), .Y(n18877) );
  NAND2X1 U12522 ( .A(n18884), .B(n18877), .Y(n18878) );
  OAI21X1 U12523 ( .A(n18879), .B(n18884), .C(n18878), .Y(n18880) );
  OAI21X1 U12524 ( .A(n18856), .B(n18891), .C(n18880), .Y(n19214) );
  INVX1 U12525 ( .A(n18881), .Y(n18883) );
  AOI22X1 U12526 ( .A(n18885), .B(n18884), .C(n18883), .D(n18882), .Y(n18894)
         );
  NAND3X1 U12527 ( .A(n18888), .B(n18887), .C(n18886), .Y(n18890) );
  AOI21X1 U12528 ( .A(n18891), .B(n18890), .C(n18889), .Y(n18892) );
  INVX1 U12529 ( .A(n18892), .Y(n18893) );
  NAND3X1 U12530 ( .A(n18895), .B(n18894), .C(n18893), .Y(n19238) );
  INVX1 U12531 ( .A(n17076), .Y(n19213) );
  AOI21X1 U12532 ( .A(n19215), .B(n16575), .C(n19213), .Y(n19206) );
  AOI21X1 U12533 ( .A(n18895), .B(n19214), .C(n19210), .Y(n19207) );
  AND2X1 U12534 ( .A(n16762), .B(n16825), .Y(n18911) );
  NAND2X1 U12535 ( .A(n18896), .B(n18944), .Y(n18931) );
  INVX1 U12536 ( .A(n18931), .Y(n18899) );
  OAI21X1 U12537 ( .A(n18899), .B(n18898), .C(n19548), .Y(n18904) );
  OAI21X1 U12538 ( .A(n16940), .B(n16473), .C(n16723), .Y(n18902) );
  INVX1 U12539 ( .A(n18902), .Y(n18909) );
  HAX1 U12540 ( .A(n18911), .B(n18908), .YS(n18903) );
  AOI22X1 U12541 ( .A(n18911), .B(n18904), .C(n18909), .D(n18903), .Y(n18914)
         );
  AOI21X1 U12542 ( .A(n16763), .B(n18905), .C(n17074), .Y(n18924) );
  AOI21X1 U12543 ( .A(n16583), .B(n18906), .C(n18924), .Y(n18907) );
  INVX1 U12544 ( .A(n18907), .Y(n18913) );
  NAND2X1 U12545 ( .A(n18909), .B(n18908), .Y(n18910) );
  AOI22X1 U12546 ( .A(n18914), .B(n18913), .C(n19342), .D(n18912), .Y(n19065)
         );
  AOI21X1 U12547 ( .A(n18784), .B(n18915), .C(n16658), .Y(n18922) );
  INVX1 U12548 ( .A(n18922), .Y(n18920) );
  NAND3X1 U12549 ( .A(n18784), .B(n19548), .C(n16512), .Y(n18918) );
  NAND3X1 U12550 ( .A(n18918), .B(n18917), .C(n16660), .Y(n18919) );
  OAI21X1 U12551 ( .A(n16660), .B(n18920), .C(n18919), .Y(n18925) );
  AOI21X1 U12552 ( .A(n16762), .B(n18922), .C(n16657), .Y(n19338) );
  INVX1 U12553 ( .A(n16428), .Y(n19332) );
  AOI22X1 U12554 ( .A(n18925), .B(n18924), .C(n17074), .D(n19332), .Y(n19064)
         );
  AND2X1 U12555 ( .A(n18927), .B(n18926), .Y(n18948) );
  NAND2X1 U12556 ( .A(n18927), .B(n18943), .Y(n18939) );
  INVX1 U12557 ( .A(n18939), .Y(n18946) );
  AOI21X1 U12558 ( .A(n18943), .B(n16379), .C(n18946), .Y(n18933) );
  NAND3X1 U12559 ( .A(n16927), .B(n18929), .C(n16735), .Y(n18930) );
  OAI21X1 U12560 ( .A(n18948), .B(n18931), .C(n18930), .Y(n18936) );
  AOI21X1 U12561 ( .A(n18934), .B(n16927), .C(n18932), .Y(n19329) );
  NAND3X1 U12562 ( .A(n19329), .B(n17096), .C(n16584), .Y(n18935) );
  OAI21X1 U12563 ( .A(n16584), .B(n18936), .C(n18935), .Y(n19046) );
  OR2X1 U12564 ( .A(n16666), .B(n19046), .Y(n19048) );
  NAND2X1 U12565 ( .A(n17077), .B(n19048), .Y(n19051) );
  NAND3X1 U12566 ( .A(n18940), .B(n18939), .C(n18938), .Y(n18942) );
  NAND2X1 U12567 ( .A(n18942), .B(n17073), .Y(n18955) );
  NAND2X1 U12568 ( .A(n16735), .B(n16625), .Y(n18947) );
  AOI22X1 U12569 ( .A(n18948), .B(n18947), .C(n18946), .D(n16658), .Y(n18951)
         );
  AND2X1 U12570 ( .A(n18952), .B(n18949), .Y(n18950) );
  AOI22X1 U12571 ( .A(n18955), .B(n17107), .C(n18951), .D(n18950), .Y(n18960)
         );
  OAI21X1 U12572 ( .A(n18955), .B(n16763), .C(n16449), .Y(n18956) );
  INVX1 U12573 ( .A(n18956), .Y(n19328) );
  NAND3X1 U12574 ( .A(n19328), .B(n18957), .C(n19523), .Y(n18958) );
  OAI21X1 U12575 ( .A(n18960), .B(n16952), .C(n18958), .Y(n19050) );
  NAND2X1 U12576 ( .A(n19048), .B(n19050), .Y(n19044) );
  NAND2X1 U12577 ( .A(n19051), .B(n19044), .Y(n19042) );
  NAND2X1 U12578 ( .A(\add_x_42/n1 ), .B(
        \lamb/scale_ts3/genblk1[2].mult/added[4] ), .Y(n18961) );
  INVX1 U12579 ( .A(\lamb/scale_ts3/genblk1[2].mult/added[3] ), .Y(n18962) );
  OR2X1 U12580 ( .A(\add_x_42/n1 ), .B(
        \lamb/scale_ts3/genblk1[2].mult/added[4] ), .Y(n18969) );
  NAND3X1 U12581 ( .A(n18961), .B(n18962), .C(n18969), .Y(n19033) );
  INVX1 U12582 ( .A(n18969), .Y(n18963) );
  NOR2X1 U12583 ( .A(n18962), .B(n18963), .Y(n18964) );
  OAI21X1 U12584 ( .A(n18964), .B(\lamb/scale_ts3/genblk1[2].mult/added[2] ), 
        .C(n16434), .Y(n18965) );
  NAND2X1 U12585 ( .A(n17053), .B(n18965), .Y(n18967) );
  MUX2X1 U12586 ( .B(\lamb/scale_ts3/genblk1[2].mult/added[4] ), .A(
        \lamb/scale_ts3/genblk1[2].mult/added[3] ), .S(\add_x_42/n1 ), .Y(
        n18966) );
  OAI21X1 U12587 ( .A(\lamb/scale_ts3/genblk1[2].mult/added[3] ), .B(
        \lamb/scale_ts3/genblk1[2].mult/added[4] ), .C(n18966), .Y(n19007) );
  INVX1 U12588 ( .A(n19007), .Y(n19031) );
  AOI22X1 U12589 ( .A(\lamb/scale_ts3/genblk1[2].mult/added[1] ), .B(n18967), 
        .C(\lamb/scale_ts3/genblk1[2].mult/added[2] ), .D(n19031), .Y(n18973)
         );
  NAND3X1 U12590 ( .A(\add_x_42/n1 ), .B(
        \lamb/scale_ts3/genblk1[2].mult/added[4] ), .C(
        \lamb/scale_ts3/genblk1[2].mult/added[3] ), .Y(n19028) );
  INVX1 U12591 ( .A(n16662), .Y(n18968) );
  NAND3X1 U12592 ( .A(\lamb/scale_ts3/genblk1[2].mult/added[3] ), .B(n16964), 
        .C(n18969), .Y(n18999) );
  INVX1 U12593 ( .A(n18970), .Y(n19094) );
  AOI21X1 U12594 ( .A(n16368), .B(n16373), .C(n19094), .Y(n19009) );
  INVX1 U12595 ( .A(n19009), .Y(n19034) );
  AOI21X1 U12596 ( .A(n18973), .B(n18999), .C(n19034), .Y(n18988) );
  INVX1 U12597 ( .A(\lamb/scale_ds3/genblk1[2].mult/added[1] ), .Y(n18993) );
  OR2X1 U12598 ( .A(\lamb/scale_ds3/genblk1[2].mult/added[4] ), .B(
        \add_x_46/n1 ), .Y(n18978) );
  NAND2X1 U12599 ( .A(\lamb/scale_ds3/genblk1[2].mult/added[3] ), .B(n18978), 
        .Y(n18974) );
  NOR2X1 U12600 ( .A(\lamb/scale_ds3/genblk1[2].mult/added[3] ), .B(n19020), 
        .Y(n18979) );
  INVX1 U12601 ( .A(n18979), .Y(n18975) );
  INVX1 U12602 ( .A(n18974), .Y(n18981) );
  NAND3X1 U12603 ( .A(\lamb/scale_ds3/genblk1[2].mult/added[1] ), .B(n18975), 
        .C(\lamb/scale_ds3/genblk1[2].mult/added[2] ), .Y(n18976) );
  OAI21X1 U12604 ( .A(\lamb/scale_ds3/genblk1[2].mult/added[2] ), .B(n18981), 
        .C(n18976), .Y(n18977) );
  AOI21X1 U12605 ( .A(n18993), .B(n17014), .C(n18977), .Y(n19027) );
  INVX1 U12606 ( .A(n19027), .Y(n18983) );
  INVX1 U12607 ( .A(n16330), .Y(n18980) );
  INVX1 U12608 ( .A(\lamb/scale_ds3/genblk1[2].mult/added[2] ), .Y(n18996) );
  AOI22X1 U12609 ( .A(\lamb/scale_ds3/genblk1[2].mult/added[1] ), .B(n18980), 
        .C(n19023), .D(n16342), .Y(n18982) );
  AND2X1 U12610 ( .A(n18993), .B(n18981), .Y(n19012) );
  NAND2X1 U12611 ( .A(n19012), .B(n16987), .Y(n18989) );
  NAND3X1 U12612 ( .A(n18983), .B(n18982), .C(n18989), .Y(n18986) );
  NAND2X1 U12613 ( .A(n18986), .B(n17033), .Y(n18987) );
  HAX1 U12614 ( .A(n18988), .B(n18987), .YS(n19073) );
  NOR3X1 U12615 ( .A(\lamb/scale_ds3/genblk1[2].mult/added[4] ), .B(
        \add_x_46/n1 ), .C(\lamb/scale_ds3/genblk1[2].mult/added[3] ), .Y(
        n19022) );
  INVX1 U12616 ( .A(n19022), .Y(n18990) );
  NAND2X1 U12617 ( .A(n18990), .B(n18989), .Y(n18995) );
  NAND3X1 U12618 ( .A(\lamb/scale_ds3/genblk1[2].mult/added[4] ), .B(
        \add_x_46/n1 ), .C(\lamb/scale_ds3/genblk1[2].mult/added[3] ), .Y(
        n18991) );
  AOI21X1 U12619 ( .A(n16342), .B(n18991), .C(n19022), .Y(n19013) );
  NAND2X1 U12620 ( .A(n18993), .B(n16330), .Y(n18994) );
  AOI22X1 U12621 ( .A(\lamb/scale_ds3/genblk1[2].mult/added[2] ), .B(n18995), 
        .C(n16970), .D(n18994), .Y(n18997) );
  NAND3X1 U12622 ( .A(n19020), .B(\lamb/scale_ds3/genblk1[2].mult/added[3] ), 
        .C(n18996), .Y(n19015) );
  AOI21X1 U12623 ( .A(n18997), .B(n19015), .C(n19025), .Y(n19004) );
  INVX1 U12624 ( .A(n16434), .Y(n19000) );
  INVX1 U12625 ( .A(\lamb/scale_ts3/genblk1[2].mult/added[2] ), .Y(n18998) );
  AOI22X1 U12626 ( .A(n19000), .B(n18999), .C(n16662), .D(n18998), .Y(n19011)
         );
  NAND2X1 U12627 ( .A(\lamb/scale_ts3/genblk1[2].mult/added[1] ), .B(n16571), 
        .Y(n19030) );
  AOI21X1 U12628 ( .A(\lamb/scale_ts3/genblk1[2].mult/added[2] ), .B(n16662), 
        .C(n19030), .Y(n19008) );
  INVX1 U12629 ( .A(n19008), .Y(n19001) );
  OAI21X1 U12630 ( .A(\lamb/scale_ts3/genblk1[2].mult/added[1] ), .B(n17053), 
        .C(n19001), .Y(n19002) );
  OAI21X1 U12631 ( .A(n19011), .B(n19002), .C(n19009), .Y(n19003) );
  HAX1 U12632 ( .A(n19004), .B(n19003), .YS(n19039) );
  INVX1 U12633 ( .A(n19039), .Y(n19058) );
  AOI22X1 U12634 ( .A(n19008), .B(n19007), .C(n16964), .D(n16571), .Y(n19010)
         );
  OAI21X1 U12635 ( .A(n19011), .B(n19010), .C(n19009), .Y(n19018) );
  AOI22X1 U12636 ( .A(\lamb/scale_ds3/genblk1[2].mult/added[1] ), .B(n19023), 
        .C(\lamb/scale_ds3/genblk1[2].mult/added[2] ), .D(n19012), .Y(n19014)
         );
  NAND3X1 U12637 ( .A(n19015), .B(n19014), .C(n16970), .Y(n19016) );
  NAND2X1 U12638 ( .A(n19016), .B(n17033), .Y(n19017) );
  HAX1 U12639 ( .A(n19018), .B(n19017), .YS(n19052) );
  INVX1 U12640 ( .A(n19052), .Y(n19061) );
  NAND2X1 U12641 ( .A(n16987), .B(n16330), .Y(n19021) );
  AOI22X1 U12642 ( .A(\lamb/scale_ds3/genblk1[2].mult/added[1] ), .B(n19022), 
        .C(\lamb/scale_ds3/genblk1[2].mult/added[2] ), .D(n19021), .Y(n19024)
         );
  AOI22X1 U12643 ( .A(\lamb/scale_ds3/genblk1[2].mult/added[1] ), .B(
        \lamb/scale_ds3/genblk1[2].mult/added[2] ), .C(n19024), .D(n17014), 
        .Y(n19026) );
  OAI21X1 U12644 ( .A(n19027), .B(n19026), .C(n17033), .Y(n19038) );
  OAI21X1 U12645 ( .A(\lamb/scale_ts3/genblk1[2].mult/added[1] ), .B(n16662), 
        .C(n17053), .Y(n19029) );
  AOI22X1 U12646 ( .A(n19031), .B(n19030), .C(
        \lamb/scale_ts3/genblk1[2].mult/added[2] ), .D(n19029), .Y(n19036) );
  NAND3X1 U12647 ( .A(\lamb/scale_ts3/genblk1[2].mult/added[1] ), .B(n17053), 
        .C(n16434), .Y(n19035) );
  AOI21X1 U12648 ( .A(n19036), .B(n19035), .C(n19034), .Y(n19037) );
  HAX1 U12649 ( .A(n19038), .B(n19037), .YS(n19062) );
  INVX1 U12650 ( .A(n19062), .Y(n19053) );
  NAND3X1 U12651 ( .A(n19053), .B(n16637), .C(n17055), .Y(n19041) );
  NAND3X1 U12652 ( .A(n16581), .B(n19041), .C(n19040), .Y(n19333) );
  AOI21X1 U12653 ( .A(n19042), .B(n16461), .C(n16715), .Y(n19082) );
  NOR3X1 U12654 ( .A(n19052), .B(n16581), .C(n19053), .Y(n19356) );
  INVX1 U12655 ( .A(n19356), .Y(n19357) );
  AND2X1 U12656 ( .A(n19082), .B(n19357), .Y(n19180) );
  NOR2X1 U12657 ( .A(n19048), .B(n19050), .Y(n19063) );
  INVX1 U12658 ( .A(n17077), .Y(n19043) );
  AOI22X1 U12659 ( .A(n17077), .B(n19044), .C(n16666), .D(n19043), .Y(n19045)
         );
  NAND2X1 U12660 ( .A(n16666), .B(n19046), .Y(n19047) );
  OAI21X1 U12661 ( .A(n19048), .B(n17077), .C(n19047), .Y(n19049) );
  AOI21X1 U12662 ( .A(n19051), .B(n19050), .C(n19049), .Y(n19076) );
  INVX1 U12663 ( .A(n19073), .Y(n19055) );
  NAND2X1 U12664 ( .A(n19053), .B(n17055), .Y(n19057) );
  AOI21X1 U12665 ( .A(n19055), .B(n16604), .C(n19054), .Y(n19056) );
  AOI21X1 U12666 ( .A(n16331), .B(n19057), .C(n16800), .Y(n19349) );
  NAND3X1 U12667 ( .A(n19058), .B(n19073), .C(n16604), .Y(n19059) );
  AOI22X1 U12668 ( .A(n19062), .B(n19061), .C(n16331), .D(n19059), .Y(n19346)
         );
  AOI21X1 U12669 ( .A(n17077), .B(n16666), .C(n19063), .Y(n19066) );
  INVX1 U12670 ( .A(n19066), .Y(n19074) );
  FAX1 U12671 ( .A(n16713), .B(n19067), .C(n17064), .YC(n19075), .YS(n19113)
         );
  INVX1 U12672 ( .A(n16375), .Y(n19084) );
  OAI21X1 U12673 ( .A(n19073), .B(n19072), .C(n16604), .Y(n19371) );
  INVX1 U12674 ( .A(n19371), .Y(n19081) );
  AOI21X1 U12675 ( .A(n19075), .B(n19074), .C(n16375), .Y(n19078) );
  NAND2X1 U12676 ( .A(n19081), .B(n19078), .Y(n19079) );
  AND2X1 U12677 ( .A(n19084), .B(n19079), .Y(n19112) );
  NOR2X1 U12678 ( .A(n19113), .B(n19112), .Y(n19114) );
  FAX1 U12679 ( .A(n16715), .B(n16696), .C(n16717), .YC(n19067), .YS(n19120)
         );
  NOR2X1 U12680 ( .A(n19120), .B(n16931), .Y(n19085) );
  INVX1 U12681 ( .A(n19113), .Y(n19119) );
  NAND2X1 U12682 ( .A(n19112), .B(n19119), .Y(n19147) );
  INVX1 U12683 ( .A(n19120), .Y(n19148) );
  NAND3X1 U12684 ( .A(n19147), .B(n19149), .C(n17070), .Y(n19083) );
  INVX1 U12685 ( .A(n19083), .Y(n19086) );
  NAND2X1 U12686 ( .A(n19085), .B(n19084), .Y(n19110) );
  AOI22X1 U12687 ( .A(n19180), .B(n16355), .C(n19086), .D(n19110), .Y(n19109)
         );
  INVX1 U12688 ( .A(\lamb/scale_ts3/genblk1[3].mult/added[1] ), .Y(n19156) );
  INVX1 U12689 ( .A(\lamb/scale_ts3/genblk1[3].mult/added[3] ), .Y(n19128) );
  OR2X1 U12690 ( .A(n19128), .B(\add_x_41/n1 ), .Y(n19087) );
  AOI22X1 U12691 ( .A(\lamb/scale_ts3/genblk1[3].mult/added[4] ), .B(
        \lamb/scale_ts3/genblk1[3].mult/added[3] ), .C(n16329), .D(n19087), 
        .Y(n19123) );
  INVX1 U12692 ( .A(n19123), .Y(n19184) );
  NOR2X1 U12693 ( .A(n19156), .B(n19184), .Y(n19091) );
  INVX1 U12694 ( .A(\lamb/scale_ts3/genblk1[3].mult/added[2] ), .Y(n19088) );
  NAND3X1 U12695 ( .A(\lamb/scale_ts3/genblk1[3].mult/added[3] ), .B(
        \lamb/scale_ts3/genblk1[3].mult/added[4] ), .C(\add_x_41/n1 ), .Y(
        n19129) );
  NOR2X1 U12696 ( .A(\lamb/scale_ts3/genblk1[3].mult/added[4] ), .B(
        \add_x_41/n1 ), .Y(n19089) );
  AOI21X1 U12697 ( .A(\add_x_41/n1 ), .B(
        \lamb/scale_ts3/genblk1[3].mult/added[4] ), .C(n19089), .Y(n19127) );
  NOR3X1 U12698 ( .A(\lamb/scale_ts3/genblk1[3].mult/added[3] ), .B(
        \lamb/scale_ts3/genblk1[3].mult/added[4] ), .C(\add_x_41/n1 ), .Y(
        n19182) );
  INVX1 U12699 ( .A(n19182), .Y(n19092) );
  NAND3X1 U12700 ( .A(\lamb/scale_ts3/genblk1[3].mult/added[2] ), .B(n16965), 
        .C(n19092), .Y(n19090) );
  OAI21X1 U12701 ( .A(n19091), .B(n16317), .C(n19090), .Y(n19132) );
  NAND2X1 U12702 ( .A(\lamb/scale_ts3/genblk1[3].mult/added[2] ), .B(
        \lamb/scale_ts3/genblk1[3].mult/added[1] ), .Y(n19124) );
  NAND3X1 U12703 ( .A(n19092), .B(n19124), .C(n16656), .Y(n19093) );
  OAI21X1 U12704 ( .A(n16656), .B(n19156), .C(n19093), .Y(n19130) );
  AOI21X1 U12705 ( .A(n19096), .B(n16372), .C(n19094), .Y(n19186) );
  INVX1 U12706 ( .A(n16358), .Y(n19131) );
  AOI21X1 U12707 ( .A(n19132), .B(n19130), .C(n19131), .Y(n19108) );
  NAND2X1 U12708 ( .A(\add_x_45/n1 ), .B(
        \lamb/scale_ds3/genblk1[3].mult/added[4] ), .Y(n19098) );
  INVX1 U12709 ( .A(\lamb/scale_ds3/genblk1[3].mult/added[3] ), .Y(n19134) );
  OR2X1 U12710 ( .A(n19134), .B(\add_x_45/n1 ), .Y(n19097) );
  AOI22X1 U12711 ( .A(\lamb/scale_ds3/genblk1[3].mult/added[4] ), .B(
        \lamb/scale_ds3/genblk1[3].mult/added[3] ), .C(n19098), .D(n19097), 
        .Y(n19190) );
  INVX1 U12712 ( .A(\lamb/scale_ds3/genblk1[3].mult/added[2] ), .Y(n19101) );
  NAND2X1 U12713 ( .A(\lamb/scale_ds3/genblk1[3].mult/added[1] ), .B(n19101), 
        .Y(n19137) );
  INVX1 U12714 ( .A(n19137), .Y(n19103) );
  NOR2X1 U12715 ( .A(\add_x_45/n1 ), .B(
        \lamb/scale_ds3/genblk1[3].mult/added[4] ), .Y(n19099) );
  AND2X1 U12716 ( .A(\lamb/scale_ds3/genblk1[3].mult/added[2] ), .B(n16602), 
        .Y(n19168) );
  AOI21X1 U12717 ( .A(\lamb/scale_ds3/genblk1[3].mult/added[4] ), .B(
        \add_x_45/n1 ), .C(n19099), .Y(n19135) );
  NAND2X1 U12718 ( .A(n19135), .B(\lamb/scale_ds3/genblk1[3].mult/added[3] ), 
        .Y(n19136) );
  OR2X1 U12719 ( .A(\lamb/scale_ds3/genblk1[3].mult/added[1] ), .B(n19136), 
        .Y(n19172) );
  AND2X1 U12720 ( .A(\lamb/scale_ds3/genblk1[3].mult/added[4] ), .B(
        \lamb/scale_ds3/genblk1[3].mult/added[3] ), .Y(n19100) );
  AOI22X1 U12721 ( .A(n19168), .B(n19172), .C(n19101), .D(n17083), .Y(n19102)
         );
  AOI21X1 U12722 ( .A(n16606), .B(n19103), .C(n19102), .Y(n19141) );
  INVX1 U12723 ( .A(\lamb/scale_ds3/genblk1[3].mult/added[1] ), .Y(n19193) );
  NAND2X1 U12724 ( .A(\lamb/scale_ds3/genblk1[3].mult/added[2] ), .B(
        \lamb/scale_ds3/genblk1[3].mult/added[1] ), .Y(n19165) );
  NAND3X1 U12725 ( .A(n19165), .B(n16602), .C(n17083), .Y(n19104) );
  OAI21X1 U12726 ( .A(n17083), .B(n19193), .C(n19104), .Y(n19138) );
  NAND2X1 U12727 ( .A(n19106), .B(n19105), .Y(n19196) );
  INVX1 U12728 ( .A(n19196), .Y(n19139) );
  AOI21X1 U12729 ( .A(n19141), .B(n19138), .C(n19139), .Y(n19107) );
  HAX1 U12730 ( .A(n16871), .B(n19107), .YS(n19378) );
  INVX1 U12731 ( .A(n19378), .Y(n19379) );
  HAX1 U12732 ( .A(n16869), .B(n19379), .YS(n19219) );
  INVX1 U12733 ( .A(n19219), .Y(n19230) );
  OAI21X1 U12734 ( .A(n19113), .B(n19149), .C(n19110), .Y(n19111) );
  AOI21X1 U12735 ( .A(n19113), .B(n17027), .C(n19111), .Y(n19122) );
  NAND2X1 U12736 ( .A(n19113), .B(n19112), .Y(n19117) );
  OAI21X1 U12737 ( .A(n19120), .B(n19114), .C(n19117), .Y(n19115) );
  OAI21X1 U12738 ( .A(n19117), .B(n19116), .C(n19115), .Y(n19121) );
  NAND3X1 U12739 ( .A(n19120), .B(n19119), .C(n16931), .Y(n19151) );
  AOI22X1 U12740 ( .A(n19180), .B(n19122), .C(n17070), .D(n16356), .Y(n19144)
         );
  NAND2X1 U12741 ( .A(\lamb/scale_ts3/genblk1[3].mult/added[2] ), .B(n19123), 
        .Y(n19158) );
  AOI21X1 U12742 ( .A(n19128), .B(n16329), .C(n19124), .Y(n19126) );
  AOI21X1 U12743 ( .A(n19156), .B(n19158), .C(n16799), .Y(n19153) );
  NAND2X1 U12744 ( .A(n19128), .B(n19127), .Y(n19157) );
  AOI22X1 U12745 ( .A(n19154), .B(n19153), .C(n19130), .D(n16959), .Y(n19133)
         );
  AOI21X1 U12746 ( .A(n19133), .B(n19132), .C(n19131), .Y(n19143) );
  NAND2X1 U12747 ( .A(n16410), .B(n17083), .Y(n19191) );
  AOI21X1 U12748 ( .A(n19138), .B(n19191), .C(n16902), .Y(n19140) );
  AOI21X1 U12749 ( .A(n19141), .B(n19140), .C(n19139), .Y(n19142) );
  HAX1 U12750 ( .A(n19143), .B(n19142), .YS(n19363) );
  HAX1 U12751 ( .A(n19144), .B(n19363), .YS(n19145) );
  INVX1 U12752 ( .A(n19145), .Y(n19225) );
  NAND3X1 U12753 ( .A(n19148), .B(n19147), .C(n17027), .Y(n19150) );
  AOI22X1 U12754 ( .A(n19180), .B(n19177), .C(n17070), .D(n16355), .Y(n19176)
         );
  OAI21X1 U12755 ( .A(n16317), .B(n19154), .C(n19153), .Y(n19181) );
  AOI21X1 U12756 ( .A(n19158), .B(n19157), .C(n19156), .Y(n19159) );
  INVX1 U12757 ( .A(n19159), .Y(n19161) );
  NAND3X1 U12758 ( .A(n19181), .B(n19161), .C(n16965), .Y(n19162) );
  NAND2X1 U12759 ( .A(n16358), .B(n19162), .Y(n19175) );
  INVX1 U12760 ( .A(n16410), .Y(n19163) );
  AOI22X1 U12761 ( .A(\lamb/scale_ds3/genblk1[3].mult/added[2] ), .B(n16606), 
        .C(\lamb/scale_ds3/genblk1[3].mult/added[1] ), .D(n19163), .Y(n19171)
         );
  AOI22X1 U12762 ( .A(n19168), .B(n16410), .C(n19166), .D(n19165), .Y(n19169)
         );
  NOR2X1 U12763 ( .A(n16902), .B(n19169), .Y(n19189) );
  NAND3X1 U12764 ( .A(n19172), .B(n19171), .C(n19189), .Y(n19173) );
  HAX1 U12765 ( .A(n19175), .B(n16851), .YS(n19396) );
  INVX1 U12766 ( .A(n19396), .Y(n19395) );
  HAX1 U12767 ( .A(n19176), .B(n19395), .YS(n19239) );
  AOI22X1 U12768 ( .A(n19180), .B(n16356), .C(n17070), .D(n19177), .Y(n19201)
         );
  INVX1 U12769 ( .A(n19181), .Y(n19188) );
  AOI22X1 U12770 ( .A(\lamb/scale_ts3/genblk1[3].mult/added[2] ), .B(n16959), 
        .C(\lamb/scale_ts3/genblk1[3].mult/added[1] ), .D(n19182), .Y(n19185)
         );
  AOI22X1 U12771 ( .A(\lamb/scale_ts3/genblk1[3].mult/added[2] ), .B(
        \lamb/scale_ts3/genblk1[3].mult/added[1] ), .C(n19185), .D(n19184), 
        .Y(n19187) );
  OAI21X1 U12772 ( .A(n19188), .B(n19187), .C(n16358), .Y(n19200) );
  INVX1 U12773 ( .A(n19189), .Y(n19198) );
  AOI21X1 U12774 ( .A(\lamb/scale_ds3/genblk1[3].mult/added[2] ), .B(n19191), 
        .C(n16606), .Y(n19195) );
  OR2X1 U12775 ( .A(n19193), .B(n16602), .Y(n19194) );
  AOI22X1 U12776 ( .A(\lamb/scale_ds3/genblk1[3].mult/added[1] ), .B(
        \lamb/scale_ds3/genblk1[3].mult/added[2] ), .C(n19195), .D(n19194), 
        .Y(n19197) );
  OAI21X1 U12777 ( .A(n19198), .B(n19197), .C(n19196), .Y(n19199) );
  HAX1 U12778 ( .A(n19200), .B(n19199), .YS(n19389) );
  HAX1 U12779 ( .A(n19201), .B(n19389), .YS(n19229) );
  NAND2X1 U12780 ( .A(n19230), .B(n19229), .Y(n19202) );
  NOR3X1 U12781 ( .A(n19221), .B(n19239), .C(n19202), .Y(n19203) );
  AOI21X1 U12782 ( .A(n16377), .B(n16367), .C(n19203), .Y(n19251) );
  NOR2X1 U12783 ( .A(n16635), .B(n17076), .Y(n19205) );
  NOR3X1 U12784 ( .A(n16367), .B(n16377), .C(n19205), .Y(n19233) );
  OAI21X1 U12785 ( .A(n19229), .B(n16615), .C(n19239), .Y(n19208) );
  AOI22X1 U12786 ( .A(n16615), .B(n19229), .C(n19208), .D(n17005), .Y(n19245)
         );
  AOI21X1 U12787 ( .A(n19214), .B(n16607), .C(n17076), .Y(n19211) );
  OAI21X1 U12788 ( .A(n19214), .B(n16607), .C(n19211), .Y(n19212) );
  NAND2X1 U12789 ( .A(n16635), .B(n19212), .Y(n19244) );
  NAND2X1 U12790 ( .A(n19245), .B(n19244), .Y(n19243) );
  INVX1 U12791 ( .A(n19243), .Y(n19249) );
  OAI21X1 U12792 ( .A(n19214), .B(n19213), .C(n16635), .Y(n19218) );
  NAND2X1 U12793 ( .A(n19214), .B(n19213), .Y(n19217) );
  AOI21X1 U12794 ( .A(n19215), .B(n17076), .C(n16575), .Y(n19216) );
  AOI21X1 U12795 ( .A(n19218), .B(n19217), .C(n19216), .Y(n19248) );
  INVX1 U12796 ( .A(n19229), .Y(n19220) );
  INVX1 U12797 ( .A(n16494), .Y(n19224) );
  INVX1 U12798 ( .A(n19239), .Y(n19226) );
  NAND2X1 U12799 ( .A(n19226), .B(n19225), .Y(n19223) );
  OAI21X1 U12800 ( .A(n19223), .B(n19224), .C(n19220), .Y(n19222) );
  AOI22X1 U12801 ( .A(n19224), .B(n19223), .C(n19222), .D(n16371), .Y(n19247)
         );
  NAND3X1 U12802 ( .A(n19226), .B(n19225), .C(n16494), .Y(n19227) );
  AOI22X1 U12803 ( .A(n19230), .B(n19229), .C(n16371), .D(n19227), .Y(n19231)
         );
  INVX1 U12804 ( .A(n19464), .Y(n19497) );
  FAX1 U12805 ( .A(n19233), .B(n19232), .C(n16595), .YC(n19458), .YS(n19464)
         );
  AND2X1 U12806 ( .A(n16635), .B(n16607), .Y(n19237) );
  OAI21X1 U12807 ( .A(n17076), .B(n19237), .C(n16575), .Y(n19457) );
  OAI21X1 U12808 ( .A(n16615), .B(n19221), .C(n19239), .Y(n19241) );
  NOR3X1 U12809 ( .A(n19458), .B(n19457), .C(n17071), .Y(n19496) );
  NOR2X1 U12810 ( .A(n19497), .B(n19496), .Y(n19452) );
  OAI21X1 U12811 ( .A(n19245), .B(n19244), .C(n19243), .Y(n19250) );
  INVX1 U12812 ( .A(n19250), .Y(n19246) );
  INVX1 U12813 ( .A(n16500), .Y(n19506) );
  AOI21X1 U12814 ( .A(n16527), .B(n19452), .C(n19506), .Y(n19255) );
  FAX1 U12815 ( .A(n19249), .B(n16697), .C(n16594), .YC(n19232), .YS(n19504)
         );
  FAX1 U12816 ( .A(n19457), .B(n17071), .C(n19458), .YC(n19498), .YS(n19252)
         );
  INVX1 U12817 ( .A(n19498), .Y(n19451) );
  NAND2X1 U12818 ( .A(n19497), .B(n19451), .Y(n19461) );
  OAI21X1 U12819 ( .A(n19504), .B(n19252), .C(n19461), .Y(n19513) );
  INVX1 U12820 ( .A(n19252), .Y(n19453) );
  NAND2X1 U12821 ( .A(n19453), .B(n19504), .Y(n19253) );
  NAND3X1 U12822 ( .A(n19514), .B(n19451), .C(n19253), .Y(n19254) );
  OAI21X1 U12823 ( .A(n19255), .B(n19513), .C(n19254), .Y(n19640) );
  AOI21X1 U12824 ( .A(n16762), .B(n19258), .C(n16657), .Y(n19263) );
  MUX2X1 U12825 ( .B(n19265), .A(n16612), .S(n16981), .Y(n19315) );
  NAND2X1 U12826 ( .A(n19272), .B(n19273), .Y(n19288) );
  AOI22X1 U12827 ( .A(n17056), .B(n16995), .C(n19280), .D(n19271), .Y(n19289)
         );
  OR2X1 U12828 ( .A(n19273), .B(n19272), .Y(n19287) );
  OAI21X1 U12829 ( .A(n16874), .B(n16455), .C(n19287), .Y(n19274) );
  NAND3X1 U12830 ( .A(n19262), .B(n19277), .C(n16360), .Y(n19276) );
  MUX2X1 U12831 ( .B(n19280), .A(n16643), .S(n19276), .Y(n19302) );
  INVX1 U12832 ( .A(n19277), .Y(n19278) );
  AOI21X1 U12833 ( .A(n16643), .B(n16360), .C(n19278), .Y(n19281) );
  OR2X1 U12834 ( .A(n16648), .B(n19281), .Y(n19283) );
  NAND2X1 U12835 ( .A(n16648), .B(n19281), .Y(n19284) );
  NAND2X1 U12836 ( .A(n17056), .B(n19284), .Y(n19286) );
  AOI21X1 U12837 ( .A(n19284), .B(n19283), .C(n17056), .Y(n19305) );
  INVX1 U12838 ( .A(n19305), .Y(n19285) );
  OAI21X1 U12839 ( .A(n16577), .B(n19286), .C(n19285), .Y(n19299) );
  HAX1 U12840 ( .A(n19290), .B(n16455), .YS(n19309) );
  OR2X1 U12841 ( .A(n19299), .B(n19309), .Y(n19292) );
  OAI21X1 U12842 ( .A(n19302), .B(n19313), .C(n19292), .Y(n19317) );
  AND2X1 U12843 ( .A(n19309), .B(n19302), .Y(n19314) );
  NAND2X1 U12844 ( .A(n19314), .B(n19299), .Y(n19291) );
  INVX1 U12845 ( .A(n19315), .Y(n19298) );
  INVX1 U12846 ( .A(n19309), .Y(n19297) );
  NOR2X1 U12847 ( .A(n19297), .B(n19302), .Y(n19304) );
  NAND2X1 U12848 ( .A(n19304), .B(n19299), .Y(n19294) );
  NAND2X1 U12849 ( .A(n19297), .B(n19302), .Y(n19293) );
  NAND2X1 U12850 ( .A(n19298), .B(n16621), .Y(n19320) );
  NAND2X1 U12851 ( .A(n19322), .B(n19320), .Y(n19295) );
  AOI22X1 U12852 ( .A(n19315), .B(n19317), .C(n19319), .D(n19295), .Y(n19296)
         );
  NAND2X1 U12853 ( .A(n16991), .B(n19296), .Y(n19325) );
  INVX1 U12854 ( .A(n19325), .Y(n19419) );
  MUX2X1 U12855 ( .B(n19299), .A(n19298), .S(n19297), .Y(n19303) );
  MUX2X1 U12856 ( .B(n19299), .A(n19309), .S(n19315), .Y(n19300) );
  OAI21X1 U12857 ( .A(n19303), .B(n19302), .C(n16791), .Y(n19323) );
  INVX1 U12858 ( .A(n19304), .Y(n19307) );
  AOI21X1 U12859 ( .A(n19307), .B(n19315), .C(n19305), .Y(n19306) );
  OAI21X1 U12860 ( .A(n19307), .B(n19315), .C(n19306), .Y(n19308) );
  MUX2X1 U12861 ( .B(n19323), .A(n19308), .S(n19313), .Y(n19398) );
  NAND3X1 U12862 ( .A(n17056), .B(n16577), .C(n19309), .Y(n19312) );
  OAI21X1 U12863 ( .A(n19314), .B(n16621), .C(n19312), .Y(n19316) );
  MUX2X1 U12864 ( .B(n19317), .A(n19316), .S(n19315), .Y(n19417) );
  INVX1 U12865 ( .A(n19417), .Y(n19318) );
  NAND2X1 U12866 ( .A(n19318), .B(n16991), .Y(n19324) );
  OR2X1 U12867 ( .A(n19398), .B(n19324), .Y(n19399) );
  NAND2X1 U12868 ( .A(n19320), .B(n19319), .Y(n19321) );
  AOI22X1 U12869 ( .A(n19313), .B(n19323), .C(n19322), .D(n19321), .Y(n19411)
         );
  INVX1 U12870 ( .A(n19411), .Y(n19418) );
  AOI21X1 U12871 ( .A(n19418), .B(n19324), .C(n19398), .Y(n19326) );
  AOI22X1 U12872 ( .A(n19419), .B(n19399), .C(n19326), .D(n19325), .Y(n19402)
         );
  OAI21X1 U12873 ( .A(n19418), .B(n19417), .C(n16991), .Y(n19440) );
  OR2X1 U12874 ( .A(n19402), .B(n19440), .Y(n19429) );
  INVX1 U12875 ( .A(n19363), .Y(n19364) );
  NAND2X1 U12876 ( .A(n16825), .B(n19328), .Y(n19330) );
  INVX1 U12877 ( .A(n19330), .Y(n19336) );
  NAND2X1 U12878 ( .A(n16428), .B(n16651), .Y(n19331) );
  OAI21X1 U12879 ( .A(n19336), .B(n17023), .C(n19331), .Y(n19372) );
  NAND3X1 U12880 ( .A(n19336), .B(n16624), .C(n19331), .Y(n19340) );
  AOI22X1 U12881 ( .A(n19342), .B(n19332), .C(n16336), .D(n19340), .Y(n19345)
         );
  INVX1 U12882 ( .A(n16461), .Y(n19355) );
  AOI22X1 U12883 ( .A(n19336), .B(n17023), .C(n19335), .D(n16651), .Y(n19354)
         );
  NAND2X1 U12884 ( .A(n19355), .B(n19354), .Y(n19353) );
  INVX1 U12885 ( .A(n19353), .Y(n19348) );
  NAND2X1 U12886 ( .A(n19336), .B(n16624), .Y(n19337) );
  OAI21X1 U12887 ( .A(n19342), .B(n16428), .C(n19337), .Y(n19339) );
  OAI21X1 U12888 ( .A(n16336), .B(n16651), .C(n16793), .Y(n19347) );
  FAX1 U12889 ( .A(n17064), .B(n16674), .C(n19344), .YC(n19373), .YS(n19368)
         );
  INVX1 U12890 ( .A(n19368), .Y(n19380) );
  FAX1 U12891 ( .A(n19371), .B(n19372), .C(n19373), .YC(n19381), .YS(n19365)
         );
  AOI21X1 U12892 ( .A(n19365), .B(n19380), .C(n19381), .Y(n19352) );
  OR2X1 U12893 ( .A(n19373), .B(n19372), .Y(n19351) );
  FAX1 U12894 ( .A(n16717), .B(n19348), .C(n19347), .YC(n19344), .YS(n19374)
         );
  AOI21X1 U12895 ( .A(n19374), .B(n19380), .C(n19365), .Y(n19350) );
  MUX2X1 U12896 ( .B(n19352), .A(n19351), .S(n19350), .Y(n19361) );
  OAI21X1 U12897 ( .A(n19355), .B(n19354), .C(n19353), .Y(n19358) );
  NAND2X1 U12898 ( .A(n19374), .B(n19380), .Y(n19359) );
  INVX1 U12899 ( .A(n19374), .Y(n19382) );
  AOI22X1 U12900 ( .A(n19381), .B(n19359), .C(n19368), .D(n19382), .Y(n19360)
         );
  NAND3X1 U12901 ( .A(n19374), .B(n19365), .C(n19380), .Y(n19385) );
  AOI22X1 U12902 ( .A(n19361), .B(n16708), .C(n19369), .D(n16969), .Y(n19362)
         );
  MUX2X1 U12903 ( .B(n19364), .A(n19363), .S(n19362), .Y(n19413) );
  INVX1 U12904 ( .A(n19365), .Y(n19367) );
  INVX1 U12905 ( .A(n19381), .Y(n19366) );
  AOI22X1 U12906 ( .A(n19382), .B(n19367), .C(n19380), .D(n19366), .Y(n19393)
         );
  NAND2X1 U12907 ( .A(n19374), .B(n19368), .Y(n19370) );
  AOI21X1 U12908 ( .A(n19381), .B(n19370), .C(n16892), .Y(n19376) );
  NOR3X1 U12909 ( .A(n19373), .B(n19372), .C(n19371), .Y(n19384) );
  NAND2X1 U12910 ( .A(n19374), .B(n19384), .Y(n19375) );
  AOI22X1 U12911 ( .A(n16708), .B(n16938), .C(n19376), .D(n19375), .Y(n19377)
         );
  MUX2X1 U12912 ( .B(n19379), .A(n19378), .S(n19377), .Y(n19397) );
  INVX1 U12913 ( .A(n19389), .Y(n19390) );
  AOI21X1 U12914 ( .A(n19381), .B(n19380), .C(n19384), .Y(n19383) );
  MUX2X1 U12915 ( .B(n19384), .A(n19383), .S(n19382), .Y(n19386) );
  AOI22X1 U12916 ( .A(n19369), .B(n16357), .C(n16708), .D(n16969), .Y(n19388)
         );
  MUX2X1 U12917 ( .B(n19390), .A(n19389), .S(n19388), .Y(n19415) );
  NOR2X1 U12918 ( .A(n19397), .B(n19415), .Y(n19425) );
  AOI22X1 U12919 ( .A(n19369), .B(n16938), .C(n16708), .D(n16357), .Y(n19394)
         );
  MUX2X1 U12920 ( .B(n19396), .A(n19395), .S(n19394), .Y(n19437) );
  NOR3X1 U12921 ( .A(n19413), .B(n19425), .C(n19437), .Y(n19404) );
  INVX1 U12922 ( .A(n19397), .Y(n19412) );
  OR2X1 U12923 ( .A(n19412), .B(n19413), .Y(n19435) );
  AND2X1 U12924 ( .A(n19435), .B(n19437), .Y(n19408) );
  OAI21X1 U12925 ( .A(n19404), .B(n19408), .C(n16929), .Y(n19428) );
  INVX1 U12926 ( .A(n19399), .Y(n19420) );
  AOI21X1 U12927 ( .A(n19418), .B(n19417), .C(n19420), .Y(n19403) );
  NAND2X1 U12928 ( .A(n19417), .B(n19398), .Y(n19409) );
  NAND2X1 U12929 ( .A(n19419), .B(n19399), .Y(n19400) );
  NAND2X1 U12930 ( .A(n16905), .B(n19400), .Y(n19401) );
  OAI21X1 U12931 ( .A(n19403), .B(n19402), .C(n19401), .Y(n19431) );
  INVX1 U12932 ( .A(n19404), .Y(n19407) );
  OR2X1 U12933 ( .A(n19437), .B(n19413), .Y(n19405) );
  OAI21X1 U12934 ( .A(n19415), .B(n19412), .C(n19405), .Y(n19406) );
  AOI22X1 U12935 ( .A(n19415), .B(n19408), .C(n19407), .D(n19406), .Y(n19430)
         );
  INVX1 U12936 ( .A(n19409), .Y(n19421) );
  AOI21X1 U12937 ( .A(n19419), .B(n16905), .C(n19420), .Y(n19441) );
  AOI21X1 U12938 ( .A(n19421), .B(n19411), .C(n19441), .Y(n19434) );
  NAND2X1 U12939 ( .A(n19413), .B(n19412), .Y(n19424) );
  INVX1 U12940 ( .A(n19424), .Y(n19416) );
  OAI21X1 U12941 ( .A(n19415), .B(n19416), .C(n19437), .Y(n19414) );
  AOI22X1 U12942 ( .A(n19416), .B(n19415), .C(n19414), .D(n19435), .Y(n19433)
         );
  NAND2X1 U12943 ( .A(n19418), .B(n19417), .Y(n19423) );
  OAI21X1 U12944 ( .A(n19421), .B(n19420), .C(n19419), .Y(n19422) );
  AND2X1 U12945 ( .A(n19423), .B(n19422), .Y(n19474) );
  NAND2X1 U12946 ( .A(n19424), .B(n19435), .Y(n19426) );
  AOI21X1 U12947 ( .A(n19437), .B(n19426), .C(n19425), .Y(n19475) );
  FAX1 U12948 ( .A(n19429), .B(n19428), .C(n19427), .YC(n19476), .YS(n19480)
         );
  NAND2X1 U12949 ( .A(n19478), .B(n19480), .Y(n19470) );
  FAX1 U12950 ( .A(n19431), .B(n16675), .C(n17008), .YC(n19427), .YS(n19489)
         );
  FAX1 U12951 ( .A(n19476), .B(n19474), .C(n17061), .YC(n19478), .YS(n19485)
         );
  NAND2X1 U12952 ( .A(n19489), .B(n19485), .Y(n19443) );
  AND2X1 U12953 ( .A(n19470), .B(n19443), .Y(n19517) );
  OAI21X1 U12954 ( .A(n19434), .B(n19433), .C(n17008), .Y(n19444) );
  INVX1 U12955 ( .A(n19444), .Y(n19442) );
  INVX1 U12956 ( .A(n19435), .Y(n19438) );
  NOR3X1 U12957 ( .A(n19438), .B(n19437), .C(n16929), .Y(n19439) );
  AOI21X1 U12958 ( .A(n19441), .B(n19440), .C(n19439), .Y(n19445) );
  AND2X1 U12959 ( .A(n19442), .B(n19445), .Y(n19516) );
  INVX1 U12960 ( .A(n19478), .Y(n19469) );
  INVX1 U12961 ( .A(n19480), .Y(n19486) );
  NAND2X1 U12962 ( .A(n19445), .B(n19444), .Y(n19467) );
  AOI21X1 U12963 ( .A(n19469), .B(n16807), .C(n19467), .Y(n19447) );
  NAND2X1 U12964 ( .A(n17061), .B(n19474), .Y(n19483) );
  INVX1 U12965 ( .A(n19483), .Y(n19482) );
  INVX1 U12966 ( .A(n19489), .Y(n19479) );
  NAND3X1 U12967 ( .A(n19476), .B(n19482), .C(n19479), .Y(n19492) );
  AOI22X1 U12968 ( .A(n19517), .B(n19516), .C(n19447), .D(n16971), .Y(n19534)
         );
  INVX1 U12969 ( .A(n19448), .Y(n19594) );
  AOI22X1 U12970 ( .A(n16707), .B(n19640), .C(n17103), .D(n16633), .Y(n19449)
         );
  MUX2X1 U12971 ( .B(msg[43]), .A(n19450), .S(n19449), .Y(decoded[43]) );
  NOR2X1 U12972 ( .A(n19451), .B(n19464), .Y(n19455) );
  INVX1 U12973 ( .A(n19504), .Y(n19459) );
  NAND2X1 U12974 ( .A(n19459), .B(n19453), .Y(n19454) );
  NOR2X1 U12975 ( .A(n19498), .B(n19452), .Y(n19499) );
  NAND3X1 U12976 ( .A(n19504), .B(n19497), .C(n19453), .Y(n19460) );
  AOI22X1 U12977 ( .A(n19455), .B(n19454), .C(n19499), .D(n16913), .Y(n19466)
         );
  NAND3X1 U12978 ( .A(n19458), .B(n19457), .C(n17071), .Y(n19500) );
  OAI21X1 U12979 ( .A(n19498), .B(n19459), .C(n19500), .Y(n19463) );
  OAI21X1 U12980 ( .A(n19504), .B(n19461), .C(n16913), .Y(n19462) );
  AOI21X1 U12981 ( .A(n19464), .B(n19463), .C(n19462), .Y(n19505) );
  NAND2X1 U12982 ( .A(n19505), .B(n19514), .Y(n19465) );
  OAI21X1 U12983 ( .A(n16500), .B(n19466), .C(n19465), .Y(n19644) );
  INVX1 U12984 ( .A(n19467), .Y(n19518) );
  INVX1 U12985 ( .A(n19485), .Y(n19468) );
  NAND3X1 U12986 ( .A(n19480), .B(n19479), .C(n19468), .Y(n19493) );
  NAND2X1 U12987 ( .A(n19469), .B(n19486), .Y(n19471) );
  NAND3X1 U12988 ( .A(n19489), .B(n19471), .C(n19470), .Y(n19473) );
  INVX1 U12989 ( .A(n19471), .Y(n19490) );
  NAND2X1 U12990 ( .A(n19490), .B(n19485), .Y(n19472) );
  NAND3X1 U12991 ( .A(n19476), .B(n17061), .C(n19474), .Y(n19477) );
  AND2X1 U12992 ( .A(n19478), .B(n19477), .Y(n19491) );
  NAND2X1 U12993 ( .A(n19480), .B(n19479), .Y(n19481) );
  MUX2X1 U12994 ( .B(n19483), .A(n19482), .S(n19481), .Y(n19484) );
  AOI22X1 U12995 ( .A(n19491), .B(n19486), .C(n19485), .D(n19484), .Y(n19487)
         );
  AOI22X1 U12996 ( .A(n19518), .B(n19495), .C(n19516), .D(n19487), .Y(n19537)
         );
  AOI22X1 U12997 ( .A(n16707), .B(n19644), .C(n17103), .D(n16634), .Y(n19488)
         );
  MUX2X1 U12998 ( .B(msg[42]), .A(n19670), .S(n19488), .Y(decoded[42]) );
  OAI21X1 U12999 ( .A(n19491), .B(n19490), .C(n19489), .Y(n19494) );
  NAND3X1 U13000 ( .A(n19494), .B(n19493), .C(n16971), .Y(n19515) );
  AOI22X1 U13001 ( .A(n19518), .B(n16352), .C(n19516), .D(n19495), .Y(n19540)
         );
  AOI21X1 U13002 ( .A(n19498), .B(n19497), .C(n19496), .Y(n19503) );
  INVX1 U13003 ( .A(n19499), .Y(n19501) );
  NAND3X1 U13004 ( .A(n19501), .B(n19500), .C(n19504), .Y(n19502) );
  OAI21X1 U13005 ( .A(n19504), .B(n19503), .C(n19502), .Y(n19510) );
  NAND2X1 U13006 ( .A(n19506), .B(n19505), .Y(n19507) );
  OAI21X1 U13007 ( .A(n17011), .B(n19510), .C(n19507), .Y(n19648) );
  AOI22X1 U13008 ( .A(n17103), .B(n16614), .C(n16707), .D(n19648), .Y(n19508)
         );
  MUX2X1 U13009 ( .B(msg[41]), .A(n19509), .S(n19508), .Y(decoded[41]) );
  OR2X1 U13010 ( .A(n16500), .B(n19510), .Y(n19512) );
  OAI21X1 U13011 ( .A(n17011), .B(n19513), .C(n19512), .Y(n19652) );
  AOI22X1 U13012 ( .A(n19518), .B(n19517), .C(n19516), .D(n16352), .Y(n19542)
         );
  AOI22X1 U13013 ( .A(n16707), .B(n19652), .C(n17103), .D(n16616), .Y(n19521)
         );
  MUX2X1 U13014 ( .B(msg[40]), .A(n19522), .S(n19521), .Y(decoded[40]) );
  NOR3X1 U13015 ( .A(n17096), .B(n16752), .C(n19620), .Y(n19530) );
  INVX1 U13016 ( .A(n16536), .Y(n19624) );
  AOI22X1 U13017 ( .A(n19530), .B(n19640), .C(n16705), .D(n19624), .Y(n19524)
         );
  MUX2X1 U13018 ( .B(msg[39]), .A(n19525), .S(n19524), .Y(decoded[39]) );
  INVX1 U13019 ( .A(n16539), .Y(n19627) );
  AOI22X1 U13020 ( .A(n16705), .B(n19627), .C(n19530), .D(n19644), .Y(n19526)
         );
  MUX2X1 U13021 ( .B(msg[38]), .A(n19527), .S(n19526), .Y(decoded[38]) );
  INVX1 U13022 ( .A(n16542), .Y(n19630) );
  AOI22X1 U13023 ( .A(n16705), .B(n19630), .C(n19530), .D(n19648), .Y(n19528)
         );
  MUX2X1 U13024 ( .B(msg[37]), .A(n19529), .S(n19528), .Y(decoded[37]) );
  INVX1 U13025 ( .A(n16545), .Y(n19634) );
  AOI22X1 U13026 ( .A(n16705), .B(n19634), .C(n19530), .D(n19652), .Y(n19532)
         );
  MUX2X1 U13027 ( .B(msg[36]), .A(n19533), .S(n19532), .Y(decoded[36]) );
  NOR3X1 U13028 ( .A(n19569), .B(n16536), .C(n16736), .Y(n19641) );
  AOI22X1 U13029 ( .A(n17103), .B(n19641), .C(n16719), .D(n19640), .Y(n19535)
         );
  MUX2X1 U13030 ( .B(msg[35]), .A(n19536), .S(n19535), .Y(decoded[35]) );
  NOR3X1 U13031 ( .A(n19569), .B(n16539), .C(n16736), .Y(n19645) );
  AOI22X1 U13032 ( .A(n17103), .B(n19645), .C(n16719), .D(n19644), .Y(n19538)
         );
  MUX2X1 U13033 ( .B(msg[34]), .A(n19539), .S(n19538), .Y(decoded[34]) );
  NOR3X1 U13034 ( .A(n19569), .B(n16542), .C(n16736), .Y(n19649) );
  AOI22X1 U13035 ( .A(n19649), .B(n17103), .C(n16719), .D(n19648), .Y(n19541)
         );
  MUX2X1 U13036 ( .B(msg[33]), .A(n19669), .S(n19541), .Y(decoded[33]) );
  NOR3X1 U13037 ( .A(n19569), .B(n16545), .C(n16736), .Y(n19654) );
  AOI22X1 U13038 ( .A(n17103), .B(n19654), .C(n16719), .D(n19652), .Y(n19545)
         );
  MUX2X1 U13039 ( .B(msg[32]), .A(n19546), .S(n19545), .Y(decoded[32]) );
  AOI21X1 U13040 ( .A(n19549), .B(n19548), .C(n19547), .Y(n19591) );
  NOR3X1 U13041 ( .A(n19620), .B(n16751), .C(n16703), .Y(n19556) );
  NOR3X1 U13042 ( .A(n16737), .B(n19594), .C(n16580), .Y(n19557) );
  AOI22X1 U13043 ( .A(n19556), .B(n19640), .C(n19557), .D(n19624), .Y(n19550)
         );
  MUX2X1 U13044 ( .B(msg[31]), .A(n19551), .S(n16868), .Y(decoded[31]) );
  AOI22X1 U13045 ( .A(n19557), .B(n19627), .C(n19556), .D(n19644), .Y(n19552)
         );
  MUX2X1 U13046 ( .B(msg[30]), .A(n19553), .S(n19552), .Y(decoded[30]) );
  AOI22X1 U13047 ( .A(n19557), .B(n19630), .C(n19556), .D(n19648), .Y(n19554)
         );
  MUX2X1 U13048 ( .B(msg[29]), .A(n19555), .S(n19554), .Y(decoded[29]) );
  AOI22X1 U13049 ( .A(n19557), .B(n19634), .C(n19556), .D(n19652), .Y(n19558)
         );
  MUX2X1 U13050 ( .B(msg[28]), .A(n19559), .S(n19558), .Y(decoded[28]) );
  AOI22X1 U13051 ( .A(n19570), .B(n16633), .C(n16720), .D(n19640), .Y(n19560)
         );
  MUX2X1 U13052 ( .B(msg[27]), .A(n19561), .S(n19560), .Y(decoded[27]) );
  AOI22X1 U13053 ( .A(n19570), .B(n16634), .C(n16720), .D(n19644), .Y(n19562)
         );
  MUX2X1 U13054 ( .B(msg[26]), .A(n19563), .S(n19562), .Y(decoded[26]) );
  AOI22X1 U13055 ( .A(n19570), .B(n16614), .C(n16720), .D(n19648), .Y(n19564)
         );
  MUX2X1 U13056 ( .B(msg[25]), .A(n19565), .S(n19564), .Y(decoded[25]) );
  AOI22X1 U13057 ( .A(n19570), .B(n16616), .C(n16720), .D(n19652), .Y(n19567)
         );
  MUX2X1 U13058 ( .B(msg[24]), .A(n19568), .S(n19567), .Y(decoded[24]) );
  NOR3X1 U13059 ( .A(n16752), .B(n19620), .C(n16703), .Y(n19577) );
  NAND2X1 U13060 ( .A(n16737), .B(n19569), .Y(n19622) );
  AOI22X1 U13061 ( .A(n19577), .B(n19640), .C(n17069), .D(n19624), .Y(n19571)
         );
  MUX2X1 U13062 ( .B(msg[23]), .A(n19572), .S(n19571), .Y(decoded[23]) );
  AOI22X1 U13063 ( .A(n17069), .B(n19627), .C(n19577), .D(n19644), .Y(n19573)
         );
  MUX2X1 U13064 ( .B(msg[22]), .A(n19574), .S(n19573), .Y(decoded[22]) );
  AOI22X1 U13065 ( .A(n17069), .B(n19630), .C(n19577), .D(n19648), .Y(n19575)
         );
  MUX2X1 U13066 ( .B(msg[21]), .A(n19576), .S(n19575), .Y(decoded[21]) );
  AOI22X1 U13067 ( .A(n17069), .B(n19634), .C(n19577), .D(n19652), .Y(n19579)
         );
  MUX2X1 U13068 ( .B(msg[20]), .A(n19580), .S(n19579), .Y(decoded[20]) );
  AOI22X1 U13069 ( .A(n19570), .B(n19641), .C(n16721), .D(n19640), .Y(n19582)
         );
  MUX2X1 U13070 ( .B(msg[19]), .A(n19583), .S(n19582), .Y(decoded[19]) );
  AOI22X1 U13071 ( .A(n19570), .B(n19645), .C(n16721), .D(n19644), .Y(n19584)
         );
  MUX2X1 U13072 ( .B(msg[18]), .A(n19585), .S(n16867), .Y(decoded[18]) );
  AOI22X1 U13073 ( .A(n19570), .B(n19649), .C(n16721), .D(n19648), .Y(n19586)
         );
  MUX2X1 U13074 ( .B(msg[17]), .A(n19587), .S(n19586), .Y(decoded[17]) );
  AOI22X1 U13075 ( .A(n19570), .B(n19654), .C(n16721), .D(n19652), .Y(n19589)
         );
  MUX2X1 U13076 ( .B(msg[16]), .A(n19590), .S(n19589), .Y(decoded[16]) );
  INVX1 U13077 ( .A(n19591), .Y(n19593) );
  NOR3X1 U13078 ( .A(n19620), .B(n16751), .C(n16704), .Y(n19602) );
  NOR3X1 U13079 ( .A(n16737), .B(n19594), .C(n16579), .Y(n19603) );
  AOI22X1 U13080 ( .A(n19602), .B(n19640), .C(n19603), .D(n19624), .Y(n19596)
         );
  MUX2X1 U13081 ( .B(msg[15]), .A(n19597), .S(n19596), .Y(decoded[15]) );
  AOI22X1 U13082 ( .A(n19603), .B(n19627), .C(n19602), .D(n19644), .Y(n19598)
         );
  MUX2X1 U13083 ( .B(msg[14]), .A(n19599), .S(n19598), .Y(decoded[14]) );
  AOI22X1 U13084 ( .A(n19603), .B(n19630), .C(n19602), .D(n19648), .Y(n19600)
         );
  MUX2X1 U13085 ( .B(msg[13]), .A(n19601), .S(n19600), .Y(decoded[13]) );
  AOI22X1 U13086 ( .A(n19603), .B(n19634), .C(n19602), .D(n19652), .Y(n19604)
         );
  MUX2X1 U13087 ( .B(msg[12]), .A(n19605), .S(n19604), .Y(decoded[12]) );
  AOI22X1 U13088 ( .A(n16718), .B(n19640), .C(n19623), .D(n16633), .Y(n19608)
         );
  MUX2X1 U13089 ( .B(msg[11]), .A(n19609), .S(n19608), .Y(decoded[11]) );
  AOI22X1 U13090 ( .A(n16718), .B(n19644), .C(n19623), .D(n16634), .Y(n19611)
         );
  MUX2X1 U13091 ( .B(msg[10]), .A(n19612), .S(n19611), .Y(decoded[10]) );
  AOI22X1 U13092 ( .A(n19623), .B(n16614), .C(n16718), .D(n19648), .Y(n19614)
         );
  MUX2X1 U13093 ( .B(msg[9]), .A(n19615), .S(n19614), .Y(decoded[9]) );
  AOI22X1 U13094 ( .A(n19623), .B(n16616), .C(n16718), .D(n19652), .Y(n19618)
         );
  MUX2X1 U13095 ( .B(msg[8]), .A(n19619), .S(n19618), .Y(decoded[8]) );
  NOR3X1 U13096 ( .A(n16752), .B(n19620), .C(n16704), .Y(n19633) );
  AOI22X1 U13097 ( .A(n19633), .B(n19640), .C(n16706), .D(n19624), .Y(n19625)
         );
  MUX2X1 U13098 ( .B(msg[7]), .A(n19626), .S(n19625), .Y(decoded[7]) );
  AOI22X1 U13099 ( .A(n16706), .B(n19627), .C(n19633), .D(n19644), .Y(n19628)
         );
  MUX2X1 U13100 ( .B(msg[6]), .A(n19629), .S(n19628), .Y(decoded[6]) );
  AOI22X1 U13101 ( .A(n16706), .B(n19630), .C(n19633), .D(n19648), .Y(n19631)
         );
  MUX2X1 U13102 ( .B(msg[5]), .A(n19632), .S(n19631), .Y(decoded[5]) );
  AOI22X1 U13103 ( .A(n16706), .B(n19634), .C(n19633), .D(n19652), .Y(n19636)
         );
  MUX2X1 U13104 ( .B(msg[4]), .A(n19637), .S(n19636), .Y(decoded[4]) );
  AOI22X1 U13105 ( .A(n19623), .B(n19641), .C(n16722), .D(n19640), .Y(n19642)
         );
  MUX2X1 U13106 ( .B(msg[3]), .A(n19643), .S(n19642), .Y(decoded[3]) );
  AOI22X1 U13107 ( .A(n19623), .B(n19645), .C(n16722), .D(n19644), .Y(n19646)
         );
  MUX2X1 U13108 ( .B(msg[2]), .A(n19647), .S(n19646), .Y(decoded[2]) );
  AOI22X1 U13109 ( .A(n19623), .B(n19649), .C(n16722), .D(n19648), .Y(n19650)
         );
  MUX2X1 U13110 ( .B(msg[1]), .A(n19651), .S(n19650), .Y(decoded[1]) );
  AOI22X1 U13111 ( .A(n19623), .B(n19654), .C(n16722), .D(n19652), .Y(n19655)
         );
  MUX2X1 U13112 ( .B(msg[0]), .A(n19656), .S(n19655), .Y(decoded[0]) );
  OAI21X1 U13113 ( .A(n19730), .B(n16497), .C(n16744), .Y(n19658) );
  INVX1 U13114 ( .A(n19660), .Y(n19662) );
  OAI21X1 U13115 ( .A(n19663), .B(n19662), .C(n17006), .Y(n9913) );
  NOR2X1 U13116 ( .A(n19699), .B(n17022), .Y(n19665) );
  NOR3X1 U13117 ( .A(n16578), .B(n19666), .C(n19665), .Y(n9912) );
  AOI22X1 U13118 ( .A(msg[59]), .B(msg[33]), .C(n19669), .D(n19668), .Y(n19673) );
  AOI22X1 U13119 ( .A(msg[42]), .B(msg[44]), .C(n19671), .D(n19670), .Y(n19672) );
  FAX1 U13120 ( .A(n19674), .B(n16676), .C(n16596), .YS(n19688) );
  INVX1 U13121 ( .A(n19686), .Y(n19685) );
  MUX2X1 U13122 ( .B(n19677), .A(n19676), .S(n17049), .Y(n19678) );
  FAX1 U13123 ( .A(n19680), .B(n19679), .C(n19678), .YS(n19681) );
  FAX1 U13124 ( .A(n17037), .B(n19682), .C(n19681), .YS(n19684) );
  MUX2X1 U13125 ( .B(n19686), .A(n19685), .S(n19684), .Y(n19687) );
  FAX1 U13126 ( .A(n19689), .B(n19688), .C(n19687), .YS(n19695) );
  MUX2X1 U13127 ( .B(n19692), .A(n19691), .S(n16378), .Y(n19693) );
  FAX1 U13128 ( .A(n19696), .B(n19695), .C(n16597), .YS(n19698) );
  OAI21X1 U13129 ( .A(n19699), .B(n19698), .C(n17047), .Y(n9911) );
  AOI22X1 U13130 ( .A(n19711), .B(n19701), .C(n19700), .D(n16422), .Y(n19702)
         );
  AOI21X1 U13131 ( .A(n19703), .B(n19710), .C(n19702), .Y(
        \lamb/scale_bs2/genblk1[1].mult/added[2] ) );
  OAI21X1 U13132 ( .A(n17080), .B(n19707), .C(n16598), .Y(n9907) );
  AOI21X1 U13133 ( .A(n19712), .B(n19713), .C(n19709), .Y(n19773) );
  NAND2X1 U13134 ( .A(n19711), .B(n19710), .Y(n19716) );
  AND2X1 U13135 ( .A(n19713), .B(n19712), .Y(n19715) );
  OAI21X1 U13136 ( .A(n19719), .B(n16939), .C(n16464), .Y(n19723) );
  NAND2X1 U13137 ( .A(n19720), .B(n19721), .Y(n19722) );
  OAI21X1 U13138 ( .A(n19724), .B(n19723), .C(n19722), .Y(n9905) );
  NAND3X1 U13139 ( .A(n16745), .B(n19726), .C(n19725), .Y(n19728) );
  OAI21X1 U13140 ( .A(\lamb/scale_ls2/genblk1[2].mult/added[2] ), .B(n19733), 
        .C(n19732), .Y(n19734) );
  NAND2X1 U13141 ( .A(n19746), .B(n19740), .Y(n19741) );
  OAI21X1 U13142 ( .A(n19743), .B(n19742), .C(n19741), .Y(n16310) );
  AOI21X1 U13143 ( .A(n19746), .B(n19745), .C(n19744), .Y(n19747) );
  MUX2X1 U13144 ( .B(n19753), .A(n19752), .S(n19751), .Y(n19755) );
  OAI21X1 U13145 ( .A(n17079), .B(n19755), .C(n16653), .Y(n16305) );
  NAND2X1 U13146 ( .A(n19758), .B(n17029), .Y(n19764) );
  OR2X1 U13147 ( .A(n19759), .B(n19765), .Y(n19760) );
  MUX2X1 U13148 ( .B(n19762), .A(n17062), .S(n19760), .Y(n19763) );
  AOI21X1 U13149 ( .A(n19765), .B(n19764), .C(n19763), .Y(n16304) );
  OAI21X1 U13150 ( .A(n19770), .B(n19769), .C(n16392), .Y(n16302) );
  OAI21X1 U13151 ( .A(n19773), .B(n19772), .C(n16422), .Y(n16301) );
  AOI21X1 U13152 ( .A(n19776), .B(n19775), .C(n16407), .Y(n19781) );
  NAND3X1 U13153 ( .A(n19778), .B(n16325), .C(n19776), .Y(n19779) );
  INVX1 U13154 ( .A(n19779), .Y(n19780) );
  NOR3X1 U13155 ( .A(n19782), .B(n19781), .C(n19780), .Y(n16299) );
endmodule

